** sch_path: /home/ttuser/tt10-analog-buffer/xschem/buffer.sch
.subckt buffer VDD VSS out in
*.PININFO VDD:B VSS:B in:I out:O
XM1 outm in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM2 outm in VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=2 m=1
XM3 out outm VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=8 m=1
XM4 out outm VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=16 m=1
.ends
.end
