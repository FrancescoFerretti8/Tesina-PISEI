** sch_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate_test.sch
**.subckt pass_gate_test OUT
*.opin OUT
x1 VDD VDD net1 IN0 VSS VSS pass_gate
V2 VDD GND 1.8
V3 VSS GND 0
x2 VDD VDD net1 IN1 VSS VSS pass_gate
x3 VDD VDD net1 IN2 VSS VSS pass_gate
x4 VSS VDD net1 IN3 VSS VDD pass_gate
V5 net2 GND pwl 15n 0 15.1n 1.8 20n 1.8 20.1n 0
V4 net3 GND pwl 10n 0 10.1n 0.6 15n 0.6 15.1n 0
C1 net1 VSS 5p m=1
R1 OUT net1 500 m=1
C2 net2 VSS 5p m=1
R2 IN0 net2 500 m=1
C3 net3 VSS 5p m=1
R3 IN1 net3 500 m=1
C4 net4 VSS 5p m=1
R4 IN2 net4 500 m=1
C5 net5 VSS 5p m=1
R5 IN3 net5 500 m=1
V1 net4 GND 1.8
R6 net5 net4 500 m=1
R7 GND net5 500 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.control
tran 100p 50n
write pass_gate_test.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  pass_gate.sym # of pins=6
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sch
.subckt pass_gate Inp VDD out Ain VSS Inn
*.ipin Inp
*.ipin Inn
*.opin out
*.ipin Ain
*.ipin VDD
*.ipin VSS
XM10 out Inp Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Ain Inn out VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
