magic
tech sky130A
magscale 1 2
timestamp 1749999514
<< viali >>
rect 2508 876 2556 1044
rect 3142 -374 3182 -210
<< metal1 >>
rect 1350 1072 2452 1164
rect 442 992 642 1042
rect 1350 992 1442 1072
rect 2490 1044 3680 1060
rect 442 900 1442 992
rect 1614 1030 1682 1036
rect 1614 966 1620 1030
rect 1676 966 1682 1030
rect 1614 960 1682 966
rect 1806 1030 1874 1036
rect 1806 966 1812 1030
rect 1868 966 1874 1030
rect 1806 960 1874 966
rect 1998 1030 2066 1036
rect 1998 966 2004 1030
rect 2060 966 2066 1030
rect 1998 960 2066 966
rect 2190 1030 2258 1036
rect 2190 966 2196 1030
rect 2252 966 2258 1030
rect 2190 960 2258 966
rect 2382 1030 2450 1036
rect 2382 966 2388 1030
rect 2444 966 2450 1030
rect 2382 960 2450 966
rect 442 842 642 900
rect 1350 808 1442 900
rect 1704 922 1784 928
rect 1704 846 1710 922
rect 1778 846 1784 922
rect 1704 838 1784 846
rect 1896 922 1976 928
rect 1896 846 1902 922
rect 1970 846 1976 922
rect 1896 838 1976 846
rect 2088 922 2168 928
rect 2088 846 2094 922
rect 2162 846 2168 922
rect 2088 838 2168 846
rect 2280 922 2360 928
rect 2280 846 2286 922
rect 2354 846 2360 922
rect 2490 876 2508 1044
rect 2556 876 3680 1044
rect 2490 860 3680 876
rect 2280 838 2360 846
rect 1350 716 2310 808
rect 3183 661 3249 667
rect 1984 456 2052 462
rect 418 368 618 430
rect 1984 368 2052 388
rect 418 300 2052 368
rect 418 230 618 300
rect 1984 266 2052 300
rect 3183 381 3249 595
rect 3490 381 3690 456
rect 3183 315 3690 381
rect 1978 198 1984 266
rect 2052 198 2058 266
rect 3183 119 3249 315
rect 3490 256 3690 315
rect 717 2 2052 68
rect 3177 53 3183 119
rect 3249 53 3255 119
rect 420 -307 620 -250
rect 717 -307 783 2
rect 1984 -130 2052 2
rect 1020 -198 3020 -130
rect 3120 -210 3696 -194
rect 420 -373 783 -307
rect 960 -240 1030 -234
rect 960 -304 966 -240
rect 1022 -304 1030 -240
rect 960 -312 1030 -304
rect 1216 -240 1286 -234
rect 1216 -304 1222 -240
rect 1278 -304 1286 -240
rect 1216 -312 1286 -304
rect 1472 -240 1542 -234
rect 1472 -304 1478 -240
rect 1534 -304 1542 -240
rect 1472 -312 1542 -304
rect 1728 -240 1798 -234
rect 1728 -304 1734 -240
rect 1790 -304 1798 -240
rect 1728 -312 1798 -304
rect 1984 -240 2054 -234
rect 1984 -304 1990 -240
rect 2046 -304 2054 -240
rect 1984 -312 2054 -304
rect 2240 -240 2310 -234
rect 2240 -304 2246 -240
rect 2302 -304 2310 -240
rect 2240 -312 2310 -304
rect 2496 -240 2566 -234
rect 2496 -304 2502 -240
rect 2558 -304 2566 -240
rect 2496 -312 2566 -304
rect 2752 -240 2822 -234
rect 2752 -304 2758 -240
rect 2814 -304 2822 -240
rect 2752 -312 2822 -304
rect 3008 -240 3078 -234
rect 3008 -304 3014 -240
rect 3070 -304 3078 -240
rect 3008 -312 3078 -304
rect 420 -450 620 -373
rect 1092 -595 1158 -366
rect 1348 -595 1414 -366
rect 1604 -595 1670 -366
rect 1860 -595 1926 -366
rect 2116 -595 2182 -366
rect 2372 -595 2438 -366
rect 2628 -595 2694 -366
rect 2884 -595 2950 -366
rect 3120 -374 3142 -210
rect 3182 -374 3696 -210
rect 3120 -394 3696 -374
rect 1092 -620 2950 -595
rect 1092 -661 2949 -620
rect 1991 -763 2057 -661
rect 1991 -829 2571 -763
rect 2637 -829 2643 -763
<< via1 >>
rect 1620 966 1676 1030
rect 1812 966 1868 1030
rect 2004 966 2060 1030
rect 2196 966 2252 1030
rect 2388 966 2444 1030
rect 1710 846 1778 922
rect 1902 846 1970 922
rect 2094 846 2162 922
rect 2286 846 2354 922
rect 3183 595 3249 661
rect 1984 388 2052 456
rect 1984 198 2052 266
rect 3183 53 3249 119
rect 966 -304 1022 -240
rect 1222 -304 1278 -240
rect 1478 -304 1534 -240
rect 1734 -304 1790 -240
rect 1990 -304 2046 -240
rect 2246 -304 2302 -240
rect 2502 -304 2558 -240
rect 2758 -304 2814 -240
rect 3014 -304 3070 -240
rect 2571 -829 2637 -763
<< metal2 >>
rect 1999 1561 2069 1563
rect 3183 1561 3249 1565
rect 1999 1495 3249 1561
rect 1999 1348 2069 1495
rect 1612 1276 2452 1348
rect 1612 1030 1684 1276
rect 1612 966 1620 1030
rect 1676 966 1684 1030
rect 1612 960 1684 966
rect 1804 1030 1876 1276
rect 1804 966 1812 1030
rect 1868 966 1876 1030
rect 1804 958 1876 966
rect 1996 1255 2069 1276
rect 1996 1030 2068 1255
rect 2188 1040 2260 1276
rect 1996 966 2004 1030
rect 2060 966 2068 1030
rect 1996 960 2068 966
rect 2186 1030 2260 1040
rect 2380 1040 2452 1276
rect 2380 1030 2454 1040
rect 2186 966 2196 1030
rect 2252 966 2258 1030
rect 2186 960 2258 966
rect 2382 966 2388 1030
rect 2444 966 2454 1030
rect 2382 960 2454 966
rect 1704 922 1786 932
rect 1704 846 1710 922
rect 1778 850 1786 922
rect 1894 922 1980 928
rect 1778 846 1788 850
rect 1704 593 1788 846
rect 1894 846 1902 922
rect 1970 846 1980 922
rect 1894 593 1980 846
rect 2086 922 2172 930
rect 2086 846 2094 922
rect 2162 846 2172 922
rect 2086 593 2172 846
rect 2276 922 2362 930
rect 2276 846 2286 922
rect 2354 846 2362 922
rect 2276 593 2362 846
rect 3183 661 3249 1495
rect 3177 595 3183 661
rect 3249 595 3255 661
rect 1704 562 2362 593
rect 1705 507 2362 562
rect 1984 456 2052 507
rect 1978 388 1984 456
rect 2052 388 2058 456
rect 1984 266 2052 272
rect 1984 140 2052 198
rect 960 72 3078 140
rect 3183 119 3249 125
rect 960 -240 1028 72
rect 960 -304 966 -240
rect 1022 -304 1028 -240
rect 960 -312 1028 -304
rect 1216 -240 1284 72
rect 1216 -304 1222 -240
rect 1278 -304 1284 -240
rect 1216 -310 1284 -304
rect 1472 -240 1540 72
rect 1472 -304 1478 -240
rect 1534 -304 1540 -240
rect 1472 -310 1540 -304
rect 1728 -240 1796 72
rect 1728 -304 1734 -240
rect 1790 -304 1796 -240
rect 1728 -312 1796 -304
rect 1984 -240 2052 72
rect 1984 -304 1990 -240
rect 2046 -304 2052 -240
rect 1984 -312 2052 -304
rect 2240 -240 2308 72
rect 2240 -304 2246 -240
rect 2302 -304 2308 -240
rect 2240 -310 2308 -304
rect 2496 -240 2564 72
rect 2496 -304 2502 -240
rect 2558 -304 2564 -240
rect 2496 -312 2564 -304
rect 2752 -240 2820 72
rect 2752 -304 2758 -240
rect 2814 -304 2820 -240
rect 2752 -312 2820 -304
rect 3008 -240 3076 72
rect 3008 -304 3014 -240
rect 3070 -304 3076 -240
rect 3008 -312 3076 -304
rect 2571 -763 2637 -757
rect 3183 -763 3249 53
rect 2637 -829 3249 -763
rect 2571 -835 2637 -829
use sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z  XM2
timestamp 1749982881
transform 1 0 2029 0 1 936
box -551 -310 551 310
use sky130_fd_pr__pfet_01v8_lvt_C3R4VJ  XM3
timestamp 1749999421
transform 1 0 2021 0 1 -302
box -1191 -284 1191 284
<< labels >>
flabel metal1 418 230 618 430 0 FreeSans 256 0 0 0 Ain
port 3 nsew
flabel metal1 442 842 642 1042 0 FreeSans 256 0 0 0 nin
port 5 nsew
flabel metal1 3490 256 3690 456 0 FreeSans 256 0 0 0 uscita
port 4 nsew
rlabel metal1 3480 860 3680 1060 1 VSS
port 7 n
rlabel metal1 420 -450 620 -250 1 pin
port 8 n
rlabel metal1 3496 -394 3696 -194 1 VDD
port 9 n
<< end >>
