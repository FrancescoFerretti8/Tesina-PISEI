** sch_path: /home/ttuser/tt10-analog-buffer/xschem/testbench.sch
**.subckt testbench out
*.opin out
x1 VDD VSS net1 in buffer
V1 VSS GND 0
V2 VDD GND 1.8
V3 in GND pwl 0 0 10n 0 10.1n 1.8 20n 1.8 20.1n 0
C1 net1 VSS 5p m=1
R1 out net1 500 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.control
tran 100p 50n
write testbench.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  buffer.sym # of pins=4
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/buffer.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/buffer.sch
.subckt buffer VDD VSS out in
*.iopin VDD
*.iopin VSS
*.ipin in
*.opin out
XM1 outm in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outm in VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 out outm VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 out outm VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
