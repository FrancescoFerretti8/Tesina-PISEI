magic
tech sky130A
magscale 1 2
timestamp 1749971960
<< error_p >>
rect -479 145 -417 151
rect -351 145 -289 151
rect -223 145 -161 151
rect -95 145 -33 151
rect 33 145 95 151
rect 161 145 223 151
rect 289 145 351 151
rect 417 145 479 151
rect -479 111 -467 145
rect -351 111 -339 145
rect -223 111 -211 145
rect -95 111 -83 145
rect 33 111 45 145
rect 161 111 173 145
rect 289 111 301 145
rect 417 111 429 145
rect -479 105 -417 111
rect -351 105 -289 111
rect -223 105 -161 111
rect -95 105 -33 111
rect 33 105 95 111
rect 161 105 223 111
rect 289 105 351 111
rect 417 105 479 111
<< nwell >>
rect -679 -284 679 284
<< pmoslvt >>
rect -483 -136 -413 64
rect -355 -136 -285 64
rect -227 -136 -157 64
rect -99 -136 -29 64
rect 29 -136 99 64
rect 157 -136 227 64
rect 285 -136 355 64
rect 413 -136 483 64
<< pdiff >>
rect -541 52 -483 64
rect -541 -124 -529 52
rect -495 -124 -483 52
rect -541 -136 -483 -124
rect -413 52 -355 64
rect -413 -124 -401 52
rect -367 -124 -355 52
rect -413 -136 -355 -124
rect -285 52 -227 64
rect -285 -124 -273 52
rect -239 -124 -227 52
rect -285 -136 -227 -124
rect -157 52 -99 64
rect -157 -124 -145 52
rect -111 -124 -99 52
rect -157 -136 -99 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 99 52 157 64
rect 99 -124 111 52
rect 145 -124 157 52
rect 99 -136 157 -124
rect 227 52 285 64
rect 227 -124 239 52
rect 273 -124 285 52
rect 227 -136 285 -124
rect 355 52 413 64
rect 355 -124 367 52
rect 401 -124 413 52
rect 355 -136 413 -124
rect 483 52 541 64
rect 483 -124 495 52
rect 529 -124 541 52
rect 483 -136 541 -124
<< pdiffc >>
rect -529 -124 -495 52
rect -401 -124 -367 52
rect -273 -124 -239 52
rect -145 -124 -111 52
rect -17 -124 17 52
rect 111 -124 145 52
rect 239 -124 273 52
rect 367 -124 401 52
rect 495 -124 529 52
<< nsubdiff >>
rect -643 214 -547 248
rect 547 214 643 248
rect -643 151 -609 214
rect 609 151 643 214
rect -643 -214 -609 -151
rect 609 -214 643 -151
rect -643 -248 -547 -214
rect 547 -248 643 -214
<< nsubdiffcont >>
rect -547 214 547 248
rect -643 -151 -609 151
rect 609 -151 643 151
rect -547 -248 547 -214
<< poly >>
rect -483 145 -413 161
rect -483 111 -467 145
rect -429 111 -413 145
rect -483 64 -413 111
rect -355 145 -285 161
rect -355 111 -339 145
rect -301 111 -285 145
rect -355 64 -285 111
rect -227 145 -157 161
rect -227 111 -211 145
rect -173 111 -157 145
rect -227 64 -157 111
rect -99 145 -29 161
rect -99 111 -83 145
rect -45 111 -29 145
rect -99 64 -29 111
rect 29 145 99 161
rect 29 111 45 145
rect 83 111 99 145
rect 29 64 99 111
rect 157 145 227 161
rect 157 111 173 145
rect 211 111 227 145
rect 157 64 227 111
rect 285 145 355 161
rect 285 111 301 145
rect 339 111 355 145
rect 285 64 355 111
rect 413 145 483 161
rect 413 111 429 145
rect 467 111 483 145
rect 413 64 483 111
rect -483 -162 -413 -136
rect -355 -162 -285 -136
rect -227 -162 -157 -136
rect -99 -162 -29 -136
rect 29 -162 99 -136
rect 157 -162 227 -136
rect 285 -162 355 -136
rect 413 -162 483 -136
<< polycont >>
rect -467 111 -429 145
rect -339 111 -301 145
rect -211 111 -173 145
rect -83 111 -45 145
rect 45 111 83 145
rect 173 111 211 145
rect 301 111 339 145
rect 429 111 467 145
<< locali >>
rect -643 214 -547 248
rect 547 214 643 248
rect -643 151 -609 214
rect 609 151 643 214
rect -483 111 -467 145
rect -429 111 -413 145
rect -355 111 -339 145
rect -301 111 -285 145
rect -227 111 -211 145
rect -173 111 -157 145
rect -99 111 -83 145
rect -45 111 -29 145
rect 29 111 45 145
rect 83 111 99 145
rect 157 111 173 145
rect 211 111 227 145
rect 285 111 301 145
rect 339 111 355 145
rect 413 111 429 145
rect 467 111 483 145
rect -529 52 -495 68
rect -529 -140 -495 -124
rect -401 52 -367 68
rect -401 -140 -367 -124
rect -273 52 -239 68
rect -273 -140 -239 -124
rect -145 52 -111 68
rect -145 -140 -111 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 111 52 145 68
rect 111 -140 145 -124
rect 239 52 273 68
rect 239 -140 273 -124
rect 367 52 401 68
rect 367 -140 401 -124
rect 495 52 529 68
rect 495 -140 529 -124
rect -643 -214 -609 -151
rect 609 -214 643 -151
rect -643 -248 -547 -214
rect 547 -248 643 -214
<< viali >>
rect -467 111 -429 145
rect -339 111 -301 145
rect -211 111 -173 145
rect -83 111 -45 145
rect 45 111 83 145
rect 173 111 211 145
rect 301 111 339 145
rect 429 111 467 145
rect -529 -124 -495 52
rect -401 -124 -367 52
rect -273 -124 -239 52
rect -145 -124 -111 52
rect -17 -124 17 52
rect 111 -124 145 52
rect 239 -124 273 52
rect 367 -124 401 52
rect 495 -124 529 52
<< metal1 >>
rect -479 145 -417 151
rect -479 111 -467 145
rect -429 111 -417 145
rect -479 105 -417 111
rect -351 145 -289 151
rect -351 111 -339 145
rect -301 111 -289 145
rect -351 105 -289 111
rect -223 145 -161 151
rect -223 111 -211 145
rect -173 111 -161 145
rect -223 105 -161 111
rect -95 145 -33 151
rect -95 111 -83 145
rect -45 111 -33 145
rect -95 105 -33 111
rect 33 145 95 151
rect 33 111 45 145
rect 83 111 95 145
rect 33 105 95 111
rect 161 145 223 151
rect 161 111 173 145
rect 211 111 223 145
rect 161 105 223 111
rect 289 145 351 151
rect 289 111 301 145
rect 339 111 351 145
rect 289 105 351 111
rect 417 145 479 151
rect 417 111 429 145
rect 467 111 479 145
rect 417 105 479 111
rect -535 52 -489 64
rect -535 -124 -529 52
rect -495 -124 -489 52
rect -535 -136 -489 -124
rect -407 52 -361 64
rect -407 -124 -401 52
rect -367 -124 -361 52
rect -407 -136 -361 -124
rect -279 52 -233 64
rect -279 -124 -273 52
rect -239 -124 -233 52
rect -279 -136 -233 -124
rect -151 52 -105 64
rect -151 -124 -145 52
rect -111 -124 -105 52
rect -151 -136 -105 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 105 52 151 64
rect 105 -124 111 52
rect 145 -124 151 52
rect 105 -136 151 -124
rect 233 52 279 64
rect 233 -124 239 52
rect 273 -124 279 52
rect 233 -136 279 -124
rect 361 52 407 64
rect 361 -124 367 52
rect 401 -124 407 52
rect 361 -136 407 -124
rect 489 52 535 64
rect 489 -124 495 52
rect 529 -124 535 52
rect 489 -136 535 -124
<< properties >>
string FIXED_BBOX -626 -231 626 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
