magic
tech sky130A
magscale 1 2
timestamp 1749999421
<< error_p >>
rect -991 145 -929 151
rect -863 145 -801 151
rect -735 145 -673 151
rect -607 145 -545 151
rect -479 145 -417 151
rect -351 145 -289 151
rect -223 145 -161 151
rect -95 145 -33 151
rect 33 145 95 151
rect 161 145 223 151
rect 289 145 351 151
rect 417 145 479 151
rect 545 145 607 151
rect 673 145 735 151
rect 801 145 863 151
rect 929 145 991 151
rect -991 111 -979 145
rect -863 111 -851 145
rect -735 111 -723 145
rect -607 111 -595 145
rect -479 111 -467 145
rect -351 111 -339 145
rect -223 111 -211 145
rect -95 111 -83 145
rect 33 111 45 145
rect 161 111 173 145
rect 289 111 301 145
rect 417 111 429 145
rect 545 111 557 145
rect 673 111 685 145
rect 801 111 813 145
rect 929 111 941 145
rect -991 105 -929 111
rect -863 105 -801 111
rect -735 105 -673 111
rect -607 105 -545 111
rect -479 105 -417 111
rect -351 105 -289 111
rect -223 105 -161 111
rect -95 105 -33 111
rect 33 105 95 111
rect 161 105 223 111
rect 289 105 351 111
rect 417 105 479 111
rect 545 105 607 111
rect 673 105 735 111
rect 801 105 863 111
rect 929 105 991 111
<< nwell >>
rect -1191 -284 1191 284
<< pmoslvt >>
rect -995 -136 -925 64
rect -867 -136 -797 64
rect -739 -136 -669 64
rect -611 -136 -541 64
rect -483 -136 -413 64
rect -355 -136 -285 64
rect -227 -136 -157 64
rect -99 -136 -29 64
rect 29 -136 99 64
rect 157 -136 227 64
rect 285 -136 355 64
rect 413 -136 483 64
rect 541 -136 611 64
rect 669 -136 739 64
rect 797 -136 867 64
rect 925 -136 995 64
<< pdiff >>
rect -1053 52 -995 64
rect -1053 -124 -1041 52
rect -1007 -124 -995 52
rect -1053 -136 -995 -124
rect -925 52 -867 64
rect -925 -124 -913 52
rect -879 -124 -867 52
rect -925 -136 -867 -124
rect -797 52 -739 64
rect -797 -124 -785 52
rect -751 -124 -739 52
rect -797 -136 -739 -124
rect -669 52 -611 64
rect -669 -124 -657 52
rect -623 -124 -611 52
rect -669 -136 -611 -124
rect -541 52 -483 64
rect -541 -124 -529 52
rect -495 -124 -483 52
rect -541 -136 -483 -124
rect -413 52 -355 64
rect -413 -124 -401 52
rect -367 -124 -355 52
rect -413 -136 -355 -124
rect -285 52 -227 64
rect -285 -124 -273 52
rect -239 -124 -227 52
rect -285 -136 -227 -124
rect -157 52 -99 64
rect -157 -124 -145 52
rect -111 -124 -99 52
rect -157 -136 -99 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 99 52 157 64
rect 99 -124 111 52
rect 145 -124 157 52
rect 99 -136 157 -124
rect 227 52 285 64
rect 227 -124 239 52
rect 273 -124 285 52
rect 227 -136 285 -124
rect 355 52 413 64
rect 355 -124 367 52
rect 401 -124 413 52
rect 355 -136 413 -124
rect 483 52 541 64
rect 483 -124 495 52
rect 529 -124 541 52
rect 483 -136 541 -124
rect 611 52 669 64
rect 611 -124 623 52
rect 657 -124 669 52
rect 611 -136 669 -124
rect 739 52 797 64
rect 739 -124 751 52
rect 785 -124 797 52
rect 739 -136 797 -124
rect 867 52 925 64
rect 867 -124 879 52
rect 913 -124 925 52
rect 867 -136 925 -124
rect 995 52 1053 64
rect 995 -124 1007 52
rect 1041 -124 1053 52
rect 995 -136 1053 -124
<< pdiffc >>
rect -1041 -124 -1007 52
rect -913 -124 -879 52
rect -785 -124 -751 52
rect -657 -124 -623 52
rect -529 -124 -495 52
rect -401 -124 -367 52
rect -273 -124 -239 52
rect -145 -124 -111 52
rect -17 -124 17 52
rect 111 -124 145 52
rect 239 -124 273 52
rect 367 -124 401 52
rect 495 -124 529 52
rect 623 -124 657 52
rect 751 -124 785 52
rect 879 -124 913 52
rect 1007 -124 1041 52
<< nsubdiff >>
rect -1155 214 -1059 248
rect 1059 214 1155 248
rect -1155 151 -1121 214
rect 1121 151 1155 214
rect -1155 -214 -1121 -151
rect 1121 -214 1155 -151
rect -1155 -248 -1059 -214
rect 1059 -248 1155 -214
<< nsubdiffcont >>
rect -1059 214 1059 248
rect -1155 -151 -1121 151
rect 1121 -151 1155 151
rect -1059 -248 1059 -214
<< poly >>
rect -995 145 -925 161
rect -995 111 -979 145
rect -941 111 -925 145
rect -995 64 -925 111
rect -867 145 -797 161
rect -867 111 -851 145
rect -813 111 -797 145
rect -867 64 -797 111
rect -739 145 -669 161
rect -739 111 -723 145
rect -685 111 -669 145
rect -739 64 -669 111
rect -611 145 -541 161
rect -611 111 -595 145
rect -557 111 -541 145
rect -611 64 -541 111
rect -483 145 -413 161
rect -483 111 -467 145
rect -429 111 -413 145
rect -483 64 -413 111
rect -355 145 -285 161
rect -355 111 -339 145
rect -301 111 -285 145
rect -355 64 -285 111
rect -227 145 -157 161
rect -227 111 -211 145
rect -173 111 -157 145
rect -227 64 -157 111
rect -99 145 -29 161
rect -99 111 -83 145
rect -45 111 -29 145
rect -99 64 -29 111
rect 29 145 99 161
rect 29 111 45 145
rect 83 111 99 145
rect 29 64 99 111
rect 157 145 227 161
rect 157 111 173 145
rect 211 111 227 145
rect 157 64 227 111
rect 285 145 355 161
rect 285 111 301 145
rect 339 111 355 145
rect 285 64 355 111
rect 413 145 483 161
rect 413 111 429 145
rect 467 111 483 145
rect 413 64 483 111
rect 541 145 611 161
rect 541 111 557 145
rect 595 111 611 145
rect 541 64 611 111
rect 669 145 739 161
rect 669 111 685 145
rect 723 111 739 145
rect 669 64 739 111
rect 797 145 867 161
rect 797 111 813 145
rect 851 111 867 145
rect 797 64 867 111
rect 925 145 995 161
rect 925 111 941 145
rect 979 111 995 145
rect 925 64 995 111
rect -995 -162 -925 -136
rect -867 -162 -797 -136
rect -739 -162 -669 -136
rect -611 -162 -541 -136
rect -483 -162 -413 -136
rect -355 -162 -285 -136
rect -227 -162 -157 -136
rect -99 -162 -29 -136
rect 29 -162 99 -136
rect 157 -162 227 -136
rect 285 -162 355 -136
rect 413 -162 483 -136
rect 541 -162 611 -136
rect 669 -162 739 -136
rect 797 -162 867 -136
rect 925 -162 995 -136
<< polycont >>
rect -979 111 -941 145
rect -851 111 -813 145
rect -723 111 -685 145
rect -595 111 -557 145
rect -467 111 -429 145
rect -339 111 -301 145
rect -211 111 -173 145
rect -83 111 -45 145
rect 45 111 83 145
rect 173 111 211 145
rect 301 111 339 145
rect 429 111 467 145
rect 557 111 595 145
rect 685 111 723 145
rect 813 111 851 145
rect 941 111 979 145
<< locali >>
rect -1155 214 -1059 248
rect 1059 214 1155 248
rect -1155 151 -1121 214
rect 1121 151 1155 214
rect -995 111 -979 145
rect -941 111 -925 145
rect -867 111 -851 145
rect -813 111 -797 145
rect -739 111 -723 145
rect -685 111 -669 145
rect -611 111 -595 145
rect -557 111 -541 145
rect -483 111 -467 145
rect -429 111 -413 145
rect -355 111 -339 145
rect -301 111 -285 145
rect -227 111 -211 145
rect -173 111 -157 145
rect -99 111 -83 145
rect -45 111 -29 145
rect 29 111 45 145
rect 83 111 99 145
rect 157 111 173 145
rect 211 111 227 145
rect 285 111 301 145
rect 339 111 355 145
rect 413 111 429 145
rect 467 111 483 145
rect 541 111 557 145
rect 595 111 611 145
rect 669 111 685 145
rect 723 111 739 145
rect 797 111 813 145
rect 851 111 867 145
rect 925 111 941 145
rect 979 111 995 145
rect -1041 52 -1007 68
rect -1041 -140 -1007 -124
rect -913 52 -879 68
rect -913 -140 -879 -124
rect -785 52 -751 68
rect -785 -140 -751 -124
rect -657 52 -623 68
rect -657 -140 -623 -124
rect -529 52 -495 68
rect -529 -140 -495 -124
rect -401 52 -367 68
rect -401 -140 -367 -124
rect -273 52 -239 68
rect -273 -140 -239 -124
rect -145 52 -111 68
rect -145 -140 -111 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 111 52 145 68
rect 111 -140 145 -124
rect 239 52 273 68
rect 239 -140 273 -124
rect 367 52 401 68
rect 367 -140 401 -124
rect 495 52 529 68
rect 495 -140 529 -124
rect 623 52 657 68
rect 623 -140 657 -124
rect 751 52 785 68
rect 751 -140 785 -124
rect 879 52 913 68
rect 879 -140 913 -124
rect 1007 52 1041 68
rect 1007 -140 1041 -124
rect -1155 -214 -1121 -151
rect 1121 -214 1155 -151
rect -1155 -248 -1059 -214
rect 1059 -248 1155 -214
<< viali >>
rect -979 111 -941 145
rect -851 111 -813 145
rect -723 111 -685 145
rect -595 111 -557 145
rect -467 111 -429 145
rect -339 111 -301 145
rect -211 111 -173 145
rect -83 111 -45 145
rect 45 111 83 145
rect 173 111 211 145
rect 301 111 339 145
rect 429 111 467 145
rect 557 111 595 145
rect 685 111 723 145
rect 813 111 851 145
rect 941 111 979 145
rect -1041 -124 -1007 52
rect -913 -124 -879 52
rect -785 -124 -751 52
rect -657 -124 -623 52
rect -529 -124 -495 52
rect -401 -124 -367 52
rect -273 -124 -239 52
rect -145 -124 -111 52
rect -17 -124 17 52
rect 111 -124 145 52
rect 239 -124 273 52
rect 367 -124 401 52
rect 495 -124 529 52
rect 623 -124 657 52
rect 751 -124 785 52
rect 879 -124 913 52
rect 1007 -124 1041 52
<< metal1 >>
rect -991 145 -929 151
rect -991 111 -979 145
rect -941 111 -929 145
rect -991 105 -929 111
rect -863 145 -801 151
rect -863 111 -851 145
rect -813 111 -801 145
rect -863 105 -801 111
rect -735 145 -673 151
rect -735 111 -723 145
rect -685 111 -673 145
rect -735 105 -673 111
rect -607 145 -545 151
rect -607 111 -595 145
rect -557 111 -545 145
rect -607 105 -545 111
rect -479 145 -417 151
rect -479 111 -467 145
rect -429 111 -417 145
rect -479 105 -417 111
rect -351 145 -289 151
rect -351 111 -339 145
rect -301 111 -289 145
rect -351 105 -289 111
rect -223 145 -161 151
rect -223 111 -211 145
rect -173 111 -161 145
rect -223 105 -161 111
rect -95 145 -33 151
rect -95 111 -83 145
rect -45 111 -33 145
rect -95 105 -33 111
rect 33 145 95 151
rect 33 111 45 145
rect 83 111 95 145
rect 33 105 95 111
rect 161 145 223 151
rect 161 111 173 145
rect 211 111 223 145
rect 161 105 223 111
rect 289 145 351 151
rect 289 111 301 145
rect 339 111 351 145
rect 289 105 351 111
rect 417 145 479 151
rect 417 111 429 145
rect 467 111 479 145
rect 417 105 479 111
rect 545 145 607 151
rect 545 111 557 145
rect 595 111 607 145
rect 545 105 607 111
rect 673 145 735 151
rect 673 111 685 145
rect 723 111 735 145
rect 673 105 735 111
rect 801 145 863 151
rect 801 111 813 145
rect 851 111 863 145
rect 801 105 863 111
rect 929 145 991 151
rect 929 111 941 145
rect 979 111 991 145
rect 929 105 991 111
rect -1047 52 -1001 64
rect -1047 -124 -1041 52
rect -1007 -124 -1001 52
rect -1047 -136 -1001 -124
rect -919 52 -873 64
rect -919 -124 -913 52
rect -879 -124 -873 52
rect -919 -136 -873 -124
rect -791 52 -745 64
rect -791 -124 -785 52
rect -751 -124 -745 52
rect -791 -136 -745 -124
rect -663 52 -617 64
rect -663 -124 -657 52
rect -623 -124 -617 52
rect -663 -136 -617 -124
rect -535 52 -489 64
rect -535 -124 -529 52
rect -495 -124 -489 52
rect -535 -136 -489 -124
rect -407 52 -361 64
rect -407 -124 -401 52
rect -367 -124 -361 52
rect -407 -136 -361 -124
rect -279 52 -233 64
rect -279 -124 -273 52
rect -239 -124 -233 52
rect -279 -136 -233 -124
rect -151 52 -105 64
rect -151 -124 -145 52
rect -111 -124 -105 52
rect -151 -136 -105 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 105 52 151 64
rect 105 -124 111 52
rect 145 -124 151 52
rect 105 -136 151 -124
rect 233 52 279 64
rect 233 -124 239 52
rect 273 -124 279 52
rect 233 -136 279 -124
rect 361 52 407 64
rect 361 -124 367 52
rect 401 -124 407 52
rect 361 -136 407 -124
rect 489 52 535 64
rect 489 -124 495 52
rect 529 -124 535 52
rect 489 -136 535 -124
rect 617 52 663 64
rect 617 -124 623 52
rect 657 -124 663 52
rect 617 -136 663 -124
rect 745 52 791 64
rect 745 -124 751 52
rect 785 -124 791 52
rect 745 -136 791 -124
rect 873 52 919 64
rect 873 -124 879 52
rect 913 -124 919 52
rect 873 -136 919 -124
rect 1001 52 1047 64
rect 1001 -124 1007 52
rect 1041 -124 1047 52
rect 1001 -136 1047 -124
<< properties >>
string FIXED_BBOX -1138 -231 1138 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
