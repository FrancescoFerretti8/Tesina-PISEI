** sch_path: /home/ttuser/tt10-analog-buffer/xschem/buffer_casa.sch
.subckt buffer_casa VDD VSS OUT IN
*.PININFO VDD:B VSS:B IN:I OUT:O
XM1 outm IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 m=1
XM2 outm IN VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM3 OUT outm VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=1 m=1
XM4 OUT outm VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 m=1
.ends
.end
