magic
tech sky130A
magscale 1 2
timestamp 1750082308
<< viali >>
rect 8493 12393 8527 12427
rect 8309 12189 8343 12223
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 8585 11713 8619 11747
rect 8217 11305 8251 11339
rect 8493 11305 8527 11339
rect 8033 11101 8067 11135
rect 7757 10761 7791 10795
rect 7941 10625 7975 10659
rect 8493 10625 8527 10659
rect 8033 10557 8067 10591
rect 8401 10421 8435 10455
rect 8033 8925 8067 8959
rect 8125 8925 8159 8959
rect 8309 8925 8343 8959
rect 8493 8857 8527 8891
rect 7849 8789 7883 8823
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 7849 6613 7883 6647
rect 8493 5253 8527 5287
rect 7941 5185 7975 5219
rect 8033 5117 8067 5151
rect 8125 5049 8159 5083
rect 7757 4981 7791 5015
rect 7665 3145 7699 3179
rect 7849 3009 7883 3043
rect 7941 2941 7975 2975
rect 8401 2941 8435 2975
rect 8125 2873 8159 2907
rect 8125 1921 8159 1955
rect 8309 1921 8343 1955
rect 8585 1853 8619 1887
rect 7757 1513 7791 1547
rect 2973 1445 3007 1479
rect 7573 1309 7607 1343
rect 2697 1241 2731 1275
<< metal1 >>
rect 1012 14714 8924 14736
rect 1012 14662 1846 14714
rect 1898 14662 1910 14714
rect 1962 14662 1974 14714
rect 2026 14662 2038 14714
rect 2090 14662 2102 14714
rect 2154 14662 3823 14714
rect 3875 14662 3887 14714
rect 3939 14662 3951 14714
rect 4003 14662 4015 14714
rect 4067 14662 4079 14714
rect 4131 14662 5800 14714
rect 5852 14662 5864 14714
rect 5916 14662 5928 14714
rect 5980 14662 5992 14714
rect 6044 14662 6056 14714
rect 6108 14662 7777 14714
rect 7829 14662 7841 14714
rect 7893 14662 7905 14714
rect 7957 14662 7969 14714
rect 8021 14662 8033 14714
rect 8085 14662 8924 14714
rect 1012 14640 8924 14662
rect 1012 14170 9079 14192
rect 1012 14118 2834 14170
rect 2886 14118 2898 14170
rect 2950 14118 2962 14170
rect 3014 14118 3026 14170
rect 3078 14118 3090 14170
rect 3142 14118 4811 14170
rect 4863 14118 4875 14170
rect 4927 14118 4939 14170
rect 4991 14118 5003 14170
rect 5055 14118 5067 14170
rect 5119 14118 6788 14170
rect 6840 14118 6852 14170
rect 6904 14118 6916 14170
rect 6968 14118 6980 14170
rect 7032 14118 7044 14170
rect 7096 14118 8765 14170
rect 8817 14118 8829 14170
rect 8881 14118 8893 14170
rect 8945 14118 8957 14170
rect 9009 14118 9021 14170
rect 9073 14118 9079 14170
rect 1012 14096 9079 14118
rect 1012 13626 8924 13648
rect 1012 13574 1846 13626
rect 1898 13574 1910 13626
rect 1962 13574 1974 13626
rect 2026 13574 2038 13626
rect 2090 13574 2102 13626
rect 2154 13574 3823 13626
rect 3875 13574 3887 13626
rect 3939 13574 3951 13626
rect 4003 13574 4015 13626
rect 4067 13574 4079 13626
rect 4131 13574 5800 13626
rect 5852 13574 5864 13626
rect 5916 13574 5928 13626
rect 5980 13574 5992 13626
rect 6044 13574 6056 13626
rect 6108 13574 7777 13626
rect 7829 13574 7841 13626
rect 7893 13574 7905 13626
rect 7957 13574 7969 13626
rect 8021 13574 8033 13626
rect 8085 13574 8924 13626
rect 1012 13552 8924 13574
rect 1012 13082 9079 13104
rect 1012 13030 2834 13082
rect 2886 13030 2898 13082
rect 2950 13030 2962 13082
rect 3014 13030 3026 13082
rect 3078 13030 3090 13082
rect 3142 13030 4811 13082
rect 4863 13030 4875 13082
rect 4927 13030 4939 13082
rect 4991 13030 5003 13082
rect 5055 13030 5067 13082
rect 5119 13030 6788 13082
rect 6840 13030 6852 13082
rect 6904 13030 6916 13082
rect 6968 13030 6980 13082
rect 7032 13030 7044 13082
rect 7096 13030 8765 13082
rect 8817 13030 8829 13082
rect 8881 13030 8893 13082
rect 8945 13030 8957 13082
rect 9009 13030 9021 13082
rect 9073 13030 9079 13082
rect 1012 13008 9079 13030
rect 1012 12538 8924 12560
rect 1012 12486 1846 12538
rect 1898 12486 1910 12538
rect 1962 12486 1974 12538
rect 2026 12486 2038 12538
rect 2090 12486 2102 12538
rect 2154 12486 3823 12538
rect 3875 12486 3887 12538
rect 3939 12486 3951 12538
rect 4003 12486 4015 12538
rect 4067 12486 4079 12538
rect 4131 12486 5800 12538
rect 5852 12486 5864 12538
rect 5916 12486 5928 12538
rect 5980 12486 5992 12538
rect 6044 12486 6056 12538
rect 6108 12486 7777 12538
rect 7829 12486 7841 12538
rect 7893 12486 7905 12538
rect 7957 12486 7969 12538
rect 8021 12486 8033 12538
rect 8085 12486 8924 12538
rect 1012 12464 8924 12486
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 8260 12396 8493 12424
rect 8260 12384 8266 12396
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8478 12220 8484 12232
rect 8343 12192 8484 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 1012 11994 9079 12016
rect 1012 11942 2834 11994
rect 2886 11942 2898 11994
rect 2950 11942 2962 11994
rect 3014 11942 3026 11994
rect 3078 11942 3090 11994
rect 3142 11942 4811 11994
rect 4863 11942 4875 11994
rect 4927 11942 4939 11994
rect 4991 11942 5003 11994
rect 5055 11942 5067 11994
rect 5119 11942 6788 11994
rect 6840 11942 6852 11994
rect 6904 11942 6916 11994
rect 6968 11942 6980 11994
rect 7032 11942 7044 11994
rect 7096 11942 8765 11994
rect 8817 11942 8829 11994
rect 8881 11942 8893 11994
rect 8945 11942 8957 11994
rect 9009 11942 9021 11994
rect 9073 11942 9079 11994
rect 1012 11920 9079 11942
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 8036 11676 8064 11707
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 8168 11716 8217 11744
rect 8168 11704 8174 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8570 11704 8576 11756
rect 8628 11704 8634 11756
rect 8386 11676 8392 11688
rect 8036 11648 8392 11676
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 1012 11450 8924 11472
rect 1012 11398 1846 11450
rect 1898 11398 1910 11450
rect 1962 11398 1974 11450
rect 2026 11398 2038 11450
rect 2090 11398 2102 11450
rect 2154 11398 3823 11450
rect 3875 11398 3887 11450
rect 3939 11398 3951 11450
rect 4003 11398 4015 11450
rect 4067 11398 4079 11450
rect 4131 11398 5800 11450
rect 5852 11398 5864 11450
rect 5916 11398 5928 11450
rect 5980 11398 5992 11450
rect 6044 11398 6056 11450
rect 6108 11398 7777 11450
rect 7829 11398 7841 11450
rect 7893 11398 7905 11450
rect 7957 11398 7969 11450
rect 8021 11398 8033 11450
rect 8085 11398 8924 11450
rect 1012 11376 8924 11398
rect 8205 11339 8263 11345
rect 8205 11305 8217 11339
rect 8251 11336 8263 11339
rect 8386 11336 8392 11348
rect 8251 11308 8392 11336
rect 8251 11305 8263 11308
rect 8205 11299 8263 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8570 11132 8576 11144
rect 8067 11104 8576 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 1012 10906 9079 10928
rect 1012 10854 2834 10906
rect 2886 10854 2898 10906
rect 2950 10854 2962 10906
rect 3014 10854 3026 10906
rect 3078 10854 3090 10906
rect 3142 10854 4811 10906
rect 4863 10854 4875 10906
rect 4927 10854 4939 10906
rect 4991 10854 5003 10906
rect 5055 10854 5067 10906
rect 5119 10854 6788 10906
rect 6840 10854 6852 10906
rect 6904 10854 6916 10906
rect 6968 10854 6980 10906
rect 7032 10854 7044 10906
rect 7096 10854 8765 10906
rect 8817 10854 8829 10906
rect 8881 10854 8893 10906
rect 8945 10854 8957 10906
rect 9009 10854 9021 10906
rect 9073 10854 9079 10906
rect 1012 10832 9079 10854
rect 7742 10752 7748 10804
rect 7800 10752 7806 10804
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 7975 10628 8064 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8036 10597 8064 10628
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 8444 10628 8493 10656
rect 8444 10616 8450 10628
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8570 10452 8576 10464
rect 8435 10424 8576 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 1012 10362 8924 10384
rect 1012 10310 1846 10362
rect 1898 10310 1910 10362
rect 1962 10310 1974 10362
rect 2026 10310 2038 10362
rect 2090 10310 2102 10362
rect 2154 10310 3823 10362
rect 3875 10310 3887 10362
rect 3939 10310 3951 10362
rect 4003 10310 4015 10362
rect 4067 10310 4079 10362
rect 4131 10310 5800 10362
rect 5852 10310 5864 10362
rect 5916 10310 5928 10362
rect 5980 10310 5992 10362
rect 6044 10310 6056 10362
rect 6108 10310 7777 10362
rect 7829 10310 7841 10362
rect 7893 10310 7905 10362
rect 7957 10310 7969 10362
rect 8021 10310 8033 10362
rect 8085 10310 8924 10362
rect 1012 10288 8924 10310
rect 1012 9818 9079 9840
rect 1012 9766 2834 9818
rect 2886 9766 2898 9818
rect 2950 9766 2962 9818
rect 3014 9766 3026 9818
rect 3078 9766 3090 9818
rect 3142 9766 4811 9818
rect 4863 9766 4875 9818
rect 4927 9766 4939 9818
rect 4991 9766 5003 9818
rect 5055 9766 5067 9818
rect 5119 9766 6788 9818
rect 6840 9766 6852 9818
rect 6904 9766 6916 9818
rect 6968 9766 6980 9818
rect 7032 9766 7044 9818
rect 7096 9766 8765 9818
rect 8817 9766 8829 9818
rect 8881 9766 8893 9818
rect 8945 9766 8957 9818
rect 9009 9766 9021 9818
rect 9073 9766 9079 9818
rect 1012 9744 9079 9766
rect 1012 9274 8924 9296
rect 1012 9222 1846 9274
rect 1898 9222 1910 9274
rect 1962 9222 1974 9274
rect 2026 9222 2038 9274
rect 2090 9222 2102 9274
rect 2154 9222 3823 9274
rect 3875 9222 3887 9274
rect 3939 9222 3951 9274
rect 4003 9222 4015 9274
rect 4067 9222 4079 9274
rect 4131 9222 5800 9274
rect 5852 9222 5864 9274
rect 5916 9222 5928 9274
rect 5980 9222 5992 9274
rect 6044 9222 6056 9274
rect 6108 9222 7777 9274
rect 7829 9222 7841 9274
rect 7893 9222 7905 9274
rect 7957 9222 7969 9274
rect 8021 9222 8033 9274
rect 8085 9222 8924 9274
rect 1012 9200 8924 9222
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 8067 8928 8125 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8386 8956 8392 8968
rect 8343 8928 8392 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 8570 8888 8576 8900
rect 8527 8860 8576 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 7834 8780 7840 8832
rect 7892 8780 7898 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8496 8820 8524 8851
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 8352 8792 8524 8820
rect 8352 8780 8358 8792
rect 1012 8730 9079 8752
rect 1012 8678 2834 8730
rect 2886 8678 2898 8730
rect 2950 8678 2962 8730
rect 3014 8678 3026 8730
rect 3078 8678 3090 8730
rect 3142 8678 4811 8730
rect 4863 8678 4875 8730
rect 4927 8678 4939 8730
rect 4991 8678 5003 8730
rect 5055 8678 5067 8730
rect 5119 8678 6788 8730
rect 6840 8678 6852 8730
rect 6904 8678 6916 8730
rect 6968 8678 6980 8730
rect 7032 8678 7044 8730
rect 7096 8678 8765 8730
rect 8817 8678 8829 8730
rect 8881 8678 8893 8730
rect 8945 8678 8957 8730
rect 9009 8678 9021 8730
rect 9073 8678 9079 8730
rect 1012 8656 9079 8678
rect 1012 8186 8924 8208
rect 1012 8134 1846 8186
rect 1898 8134 1910 8186
rect 1962 8134 1974 8186
rect 2026 8134 2038 8186
rect 2090 8134 2102 8186
rect 2154 8134 3823 8186
rect 3875 8134 3887 8186
rect 3939 8134 3951 8186
rect 4003 8134 4015 8186
rect 4067 8134 4079 8186
rect 4131 8134 5800 8186
rect 5852 8134 5864 8186
rect 5916 8134 5928 8186
rect 5980 8134 5992 8186
rect 6044 8134 6056 8186
rect 6108 8134 7777 8186
rect 7829 8134 7841 8186
rect 7893 8134 7905 8186
rect 7957 8134 7969 8186
rect 8021 8134 8033 8186
rect 8085 8134 8924 8186
rect 1012 8112 8924 8134
rect 1012 7642 9079 7664
rect 1012 7590 2834 7642
rect 2886 7590 2898 7642
rect 2950 7590 2962 7642
rect 3014 7590 3026 7642
rect 3078 7590 3090 7642
rect 3142 7590 4811 7642
rect 4863 7590 4875 7642
rect 4927 7590 4939 7642
rect 4991 7590 5003 7642
rect 5055 7590 5067 7642
rect 5119 7590 6788 7642
rect 6840 7590 6852 7642
rect 6904 7590 6916 7642
rect 6968 7590 6980 7642
rect 7032 7590 7044 7642
rect 7096 7590 8765 7642
rect 8817 7590 8829 7642
rect 8881 7590 8893 7642
rect 8945 7590 8957 7642
rect 9009 7590 9021 7642
rect 9073 7590 9079 7642
rect 1012 7568 9079 7590
rect 1012 7098 8924 7120
rect 1012 7046 1846 7098
rect 1898 7046 1910 7098
rect 1962 7046 1974 7098
rect 2026 7046 2038 7098
rect 2090 7046 2102 7098
rect 2154 7046 3823 7098
rect 3875 7046 3887 7098
rect 3939 7046 3951 7098
rect 4003 7046 4015 7098
rect 4067 7046 4079 7098
rect 4131 7046 5800 7098
rect 5852 7046 5864 7098
rect 5916 7046 5928 7098
rect 5980 7046 5992 7098
rect 6044 7046 6056 7098
rect 6108 7046 7777 7098
rect 7829 7046 7841 7098
rect 7893 7046 7905 7098
rect 7957 7046 7969 7098
rect 8021 7046 8033 7098
rect 8085 7046 8924 7098
rect 1012 7024 8924 7046
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 8067 6752 8125 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 7834 6604 7840 6656
rect 7892 6604 7898 6656
rect 1012 6554 9079 6576
rect 1012 6502 2834 6554
rect 2886 6502 2898 6554
rect 2950 6502 2962 6554
rect 3014 6502 3026 6554
rect 3078 6502 3090 6554
rect 3142 6502 4811 6554
rect 4863 6502 4875 6554
rect 4927 6502 4939 6554
rect 4991 6502 5003 6554
rect 5055 6502 5067 6554
rect 5119 6502 6788 6554
rect 6840 6502 6852 6554
rect 6904 6502 6916 6554
rect 6968 6502 6980 6554
rect 7032 6502 7044 6554
rect 7096 6502 8765 6554
rect 8817 6502 8829 6554
rect 8881 6502 8893 6554
rect 8945 6502 8957 6554
rect 9009 6502 9021 6554
rect 9073 6502 9079 6554
rect 1012 6480 9079 6502
rect 1012 6010 8924 6032
rect 1012 5958 1846 6010
rect 1898 5958 1910 6010
rect 1962 5958 1974 6010
rect 2026 5958 2038 6010
rect 2090 5958 2102 6010
rect 2154 5958 3823 6010
rect 3875 5958 3887 6010
rect 3939 5958 3951 6010
rect 4003 5958 4015 6010
rect 4067 5958 4079 6010
rect 4131 5958 5800 6010
rect 5852 5958 5864 6010
rect 5916 5958 5928 6010
rect 5980 5958 5992 6010
rect 6044 5958 6056 6010
rect 6108 5958 7777 6010
rect 7829 5958 7841 6010
rect 7893 5958 7905 6010
rect 7957 5958 7969 6010
rect 8021 5958 8033 6010
rect 8085 5958 8924 6010
rect 1012 5936 8924 5958
rect 1012 5466 9079 5488
rect 1012 5414 2834 5466
rect 2886 5414 2898 5466
rect 2950 5414 2962 5466
rect 3014 5414 3026 5466
rect 3078 5414 3090 5466
rect 3142 5414 4811 5466
rect 4863 5414 4875 5466
rect 4927 5414 4939 5466
rect 4991 5414 5003 5466
rect 5055 5414 5067 5466
rect 5119 5414 6788 5466
rect 6840 5414 6852 5466
rect 6904 5414 6916 5466
rect 6968 5414 6980 5466
rect 7032 5414 7044 5466
rect 7096 5414 8765 5466
rect 8817 5414 8829 5466
rect 8881 5414 8893 5466
rect 8945 5414 8957 5466
rect 9009 5414 9021 5466
rect 9073 5414 9079 5466
rect 1012 5392 9079 5414
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 8444 5256 8493 5284
rect 8444 5244 8450 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 8481 5247 8539 5253
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 7944 5148 7972 5179
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7944 5120 8033 5148
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8113 5083 8171 5089
rect 8113 5049 8125 5083
rect 8159 5080 8171 5083
rect 8294 5080 8300 5092
rect 8159 5052 8300 5080
rect 8159 5049 8171 5052
rect 8113 5043 8171 5049
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 8202 5012 8208 5024
rect 7791 4984 8208 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 1012 4922 8924 4944
rect 1012 4870 1846 4922
rect 1898 4870 1910 4922
rect 1962 4870 1974 4922
rect 2026 4870 2038 4922
rect 2090 4870 2102 4922
rect 2154 4870 3823 4922
rect 3875 4870 3887 4922
rect 3939 4870 3951 4922
rect 4003 4870 4015 4922
rect 4067 4870 4079 4922
rect 4131 4870 5800 4922
rect 5852 4870 5864 4922
rect 5916 4870 5928 4922
rect 5980 4870 5992 4922
rect 6044 4870 6056 4922
rect 6108 4870 7777 4922
rect 7829 4870 7841 4922
rect 7893 4870 7905 4922
rect 7957 4870 7969 4922
rect 8021 4870 8033 4922
rect 8085 4870 8924 4922
rect 1012 4848 8924 4870
rect 1012 4378 9079 4400
rect 1012 4326 2834 4378
rect 2886 4326 2898 4378
rect 2950 4326 2962 4378
rect 3014 4326 3026 4378
rect 3078 4326 3090 4378
rect 3142 4326 4811 4378
rect 4863 4326 4875 4378
rect 4927 4326 4939 4378
rect 4991 4326 5003 4378
rect 5055 4326 5067 4378
rect 5119 4326 6788 4378
rect 6840 4326 6852 4378
rect 6904 4326 6916 4378
rect 6968 4326 6980 4378
rect 7032 4326 7044 4378
rect 7096 4326 8765 4378
rect 8817 4326 8829 4378
rect 8881 4326 8893 4378
rect 8945 4326 8957 4378
rect 9009 4326 9021 4378
rect 9073 4326 9079 4378
rect 1012 4304 9079 4326
rect 1012 3834 8924 3856
rect 1012 3782 1846 3834
rect 1898 3782 1910 3834
rect 1962 3782 1974 3834
rect 2026 3782 2038 3834
rect 2090 3782 2102 3834
rect 2154 3782 3823 3834
rect 3875 3782 3887 3834
rect 3939 3782 3951 3834
rect 4003 3782 4015 3834
rect 4067 3782 4079 3834
rect 4131 3782 5800 3834
rect 5852 3782 5864 3834
rect 5916 3782 5928 3834
rect 5980 3782 5992 3834
rect 6044 3782 6056 3834
rect 6108 3782 7777 3834
rect 7829 3782 7841 3834
rect 7893 3782 7905 3834
rect 7957 3782 7969 3834
rect 8021 3782 8033 3834
rect 8085 3782 8924 3834
rect 1012 3760 8924 3782
rect 1012 3290 9079 3312
rect 1012 3238 2834 3290
rect 2886 3238 2898 3290
rect 2950 3238 2962 3290
rect 3014 3238 3026 3290
rect 3078 3238 3090 3290
rect 3142 3238 4811 3290
rect 4863 3238 4875 3290
rect 4927 3238 4939 3290
rect 4991 3238 5003 3290
rect 5055 3238 5067 3290
rect 5119 3238 6788 3290
rect 6840 3238 6852 3290
rect 6904 3238 6916 3290
rect 6968 3238 6980 3290
rect 7032 3238 7044 3290
rect 7096 3238 8765 3290
rect 8817 3238 8829 3290
rect 8881 3238 8893 3290
rect 8945 3238 8957 3290
rect 9009 3238 9021 3290
rect 9073 3238 9079 3290
rect 1012 3216 9079 3238
rect 7650 3136 7656 3188
rect 7708 3136 7714 3188
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 7883 3012 7972 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7944 2981 7972 3012
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8352 3012 8432 3040
rect 8352 3000 8358 3012
rect 8404 2981 8432 3012
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 8294 2904 8300 2916
rect 8168 2876 8300 2904
rect 8168 2864 8174 2876
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 8404 2848 8432 2935
rect 8386 2796 8392 2848
rect 8444 2796 8450 2848
rect 1012 2746 8924 2768
rect 1012 2694 1846 2746
rect 1898 2694 1910 2746
rect 1962 2694 1974 2746
rect 2026 2694 2038 2746
rect 2090 2694 2102 2746
rect 2154 2694 3823 2746
rect 3875 2694 3887 2746
rect 3939 2694 3951 2746
rect 4003 2694 4015 2746
rect 4067 2694 4079 2746
rect 4131 2694 5800 2746
rect 5852 2694 5864 2746
rect 5916 2694 5928 2746
rect 5980 2694 5992 2746
rect 6044 2694 6056 2746
rect 6108 2694 7777 2746
rect 7829 2694 7841 2746
rect 7893 2694 7905 2746
rect 7957 2694 7969 2746
rect 8021 2694 8033 2746
rect 8085 2694 8924 2746
rect 1012 2672 8924 2694
rect 1012 2202 9079 2224
rect 1012 2150 2834 2202
rect 2886 2150 2898 2202
rect 2950 2150 2962 2202
rect 3014 2150 3026 2202
rect 3078 2150 3090 2202
rect 3142 2150 4811 2202
rect 4863 2150 4875 2202
rect 4927 2150 4939 2202
rect 4991 2150 5003 2202
rect 5055 2150 5067 2202
rect 5119 2150 6788 2202
rect 6840 2150 6852 2202
rect 6904 2150 6916 2202
rect 6968 2150 6980 2202
rect 7032 2150 7044 2202
rect 7096 2150 8765 2202
rect 8817 2150 8829 2202
rect 8881 2150 8893 2202
rect 8945 2150 8957 2202
rect 9009 2150 9021 2202
rect 9073 2150 9079 2202
rect 1012 2128 9079 2150
rect 8110 1912 8116 1964
rect 8168 1912 8174 1964
rect 8294 1912 8300 1964
rect 8352 1912 8358 1964
rect 8573 1887 8631 1893
rect 8573 1853 8585 1887
rect 8619 1884 8631 1887
rect 9306 1884 9312 1896
rect 8619 1856 9312 1884
rect 8619 1853 8631 1856
rect 8573 1847 8631 1853
rect 9306 1844 9312 1856
rect 9364 1844 9370 1896
rect 1012 1658 8924 1680
rect 1012 1606 1846 1658
rect 1898 1606 1910 1658
rect 1962 1606 1974 1658
rect 2026 1606 2038 1658
rect 2090 1606 2102 1658
rect 2154 1606 3823 1658
rect 3875 1606 3887 1658
rect 3939 1606 3951 1658
rect 4003 1606 4015 1658
rect 4067 1606 4079 1658
rect 4131 1606 5800 1658
rect 5852 1606 5864 1658
rect 5916 1606 5928 1658
rect 5980 1606 5992 1658
rect 6044 1606 6056 1658
rect 6108 1606 7777 1658
rect 7829 1606 7841 1658
rect 7893 1606 7905 1658
rect 7957 1606 7969 1658
rect 8021 1606 8033 1658
rect 8085 1606 8924 1658
rect 1012 1584 8924 1606
rect 7745 1547 7803 1553
rect 7745 1513 7757 1547
rect 7791 1544 7803 1547
rect 8110 1544 8116 1556
rect 7791 1516 8116 1544
rect 7791 1513 7803 1516
rect 7745 1507 7803 1513
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 2961 1479 3019 1485
rect 2961 1445 2973 1479
rect 3007 1476 3019 1479
rect 8294 1476 8300 1488
rect 3007 1448 8300 1476
rect 3007 1445 3019 1448
rect 2961 1439 3019 1445
rect 8294 1436 8300 1448
rect 8352 1436 8358 1488
rect 7466 1300 7472 1352
rect 7524 1340 7530 1352
rect 7561 1343 7619 1349
rect 7561 1340 7573 1343
rect 7524 1312 7573 1340
rect 7524 1300 7530 1312
rect 7561 1309 7573 1312
rect 7607 1309 7619 1343
rect 7561 1303 7619 1309
rect 2498 1232 2504 1284
rect 2556 1272 2562 1284
rect 2685 1275 2743 1281
rect 2685 1272 2697 1275
rect 2556 1244 2697 1272
rect 2556 1232 2562 1244
rect 2685 1241 2697 1244
rect 2731 1241 2743 1275
rect 2685 1235 2743 1241
rect 1012 1114 9079 1136
rect 1012 1062 2834 1114
rect 2886 1062 2898 1114
rect 2950 1062 2962 1114
rect 3014 1062 3026 1114
rect 3078 1062 3090 1114
rect 3142 1062 4811 1114
rect 4863 1062 4875 1114
rect 4927 1062 4939 1114
rect 4991 1062 5003 1114
rect 5055 1062 5067 1114
rect 5119 1062 6788 1114
rect 6840 1062 6852 1114
rect 6904 1062 6916 1114
rect 6968 1062 6980 1114
rect 7032 1062 7044 1114
rect 7096 1062 8765 1114
rect 8817 1062 8829 1114
rect 8881 1062 8893 1114
rect 8945 1062 8957 1114
rect 9009 1062 9021 1114
rect 9073 1062 9079 1114
rect 1012 1040 9079 1062
<< via1 >>
rect 1846 14662 1898 14714
rect 1910 14662 1962 14714
rect 1974 14662 2026 14714
rect 2038 14662 2090 14714
rect 2102 14662 2154 14714
rect 3823 14662 3875 14714
rect 3887 14662 3939 14714
rect 3951 14662 4003 14714
rect 4015 14662 4067 14714
rect 4079 14662 4131 14714
rect 5800 14662 5852 14714
rect 5864 14662 5916 14714
rect 5928 14662 5980 14714
rect 5992 14662 6044 14714
rect 6056 14662 6108 14714
rect 7777 14662 7829 14714
rect 7841 14662 7893 14714
rect 7905 14662 7957 14714
rect 7969 14662 8021 14714
rect 8033 14662 8085 14714
rect 2834 14118 2886 14170
rect 2898 14118 2950 14170
rect 2962 14118 3014 14170
rect 3026 14118 3078 14170
rect 3090 14118 3142 14170
rect 4811 14118 4863 14170
rect 4875 14118 4927 14170
rect 4939 14118 4991 14170
rect 5003 14118 5055 14170
rect 5067 14118 5119 14170
rect 6788 14118 6840 14170
rect 6852 14118 6904 14170
rect 6916 14118 6968 14170
rect 6980 14118 7032 14170
rect 7044 14118 7096 14170
rect 8765 14118 8817 14170
rect 8829 14118 8881 14170
rect 8893 14118 8945 14170
rect 8957 14118 9009 14170
rect 9021 14118 9073 14170
rect 1846 13574 1898 13626
rect 1910 13574 1962 13626
rect 1974 13574 2026 13626
rect 2038 13574 2090 13626
rect 2102 13574 2154 13626
rect 3823 13574 3875 13626
rect 3887 13574 3939 13626
rect 3951 13574 4003 13626
rect 4015 13574 4067 13626
rect 4079 13574 4131 13626
rect 5800 13574 5852 13626
rect 5864 13574 5916 13626
rect 5928 13574 5980 13626
rect 5992 13574 6044 13626
rect 6056 13574 6108 13626
rect 7777 13574 7829 13626
rect 7841 13574 7893 13626
rect 7905 13574 7957 13626
rect 7969 13574 8021 13626
rect 8033 13574 8085 13626
rect 2834 13030 2886 13082
rect 2898 13030 2950 13082
rect 2962 13030 3014 13082
rect 3026 13030 3078 13082
rect 3090 13030 3142 13082
rect 4811 13030 4863 13082
rect 4875 13030 4927 13082
rect 4939 13030 4991 13082
rect 5003 13030 5055 13082
rect 5067 13030 5119 13082
rect 6788 13030 6840 13082
rect 6852 13030 6904 13082
rect 6916 13030 6968 13082
rect 6980 13030 7032 13082
rect 7044 13030 7096 13082
rect 8765 13030 8817 13082
rect 8829 13030 8881 13082
rect 8893 13030 8945 13082
rect 8957 13030 9009 13082
rect 9021 13030 9073 13082
rect 1846 12486 1898 12538
rect 1910 12486 1962 12538
rect 1974 12486 2026 12538
rect 2038 12486 2090 12538
rect 2102 12486 2154 12538
rect 3823 12486 3875 12538
rect 3887 12486 3939 12538
rect 3951 12486 4003 12538
rect 4015 12486 4067 12538
rect 4079 12486 4131 12538
rect 5800 12486 5852 12538
rect 5864 12486 5916 12538
rect 5928 12486 5980 12538
rect 5992 12486 6044 12538
rect 6056 12486 6108 12538
rect 7777 12486 7829 12538
rect 7841 12486 7893 12538
rect 7905 12486 7957 12538
rect 7969 12486 8021 12538
rect 8033 12486 8085 12538
rect 8208 12384 8260 12436
rect 8484 12180 8536 12232
rect 2834 11942 2886 11994
rect 2898 11942 2950 11994
rect 2962 11942 3014 11994
rect 3026 11942 3078 11994
rect 3090 11942 3142 11994
rect 4811 11942 4863 11994
rect 4875 11942 4927 11994
rect 4939 11942 4991 11994
rect 5003 11942 5055 11994
rect 5067 11942 5119 11994
rect 6788 11942 6840 11994
rect 6852 11942 6904 11994
rect 6916 11942 6968 11994
rect 6980 11942 7032 11994
rect 7044 11942 7096 11994
rect 8765 11942 8817 11994
rect 8829 11942 8881 11994
rect 8893 11942 8945 11994
rect 8957 11942 9009 11994
rect 9021 11942 9073 11994
rect 8116 11704 8168 11756
rect 8576 11747 8628 11756
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 8392 11636 8444 11688
rect 1846 11398 1898 11450
rect 1910 11398 1962 11450
rect 1974 11398 2026 11450
rect 2038 11398 2090 11450
rect 2102 11398 2154 11450
rect 3823 11398 3875 11450
rect 3887 11398 3939 11450
rect 3951 11398 4003 11450
rect 4015 11398 4067 11450
rect 4079 11398 4131 11450
rect 5800 11398 5852 11450
rect 5864 11398 5916 11450
rect 5928 11398 5980 11450
rect 5992 11398 6044 11450
rect 6056 11398 6108 11450
rect 7777 11398 7829 11450
rect 7841 11398 7893 11450
rect 7905 11398 7957 11450
rect 7969 11398 8021 11450
rect 8033 11398 8085 11450
rect 8392 11296 8444 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8576 11092 8628 11144
rect 2834 10854 2886 10906
rect 2898 10854 2950 10906
rect 2962 10854 3014 10906
rect 3026 10854 3078 10906
rect 3090 10854 3142 10906
rect 4811 10854 4863 10906
rect 4875 10854 4927 10906
rect 4939 10854 4991 10906
rect 5003 10854 5055 10906
rect 5067 10854 5119 10906
rect 6788 10854 6840 10906
rect 6852 10854 6904 10906
rect 6916 10854 6968 10906
rect 6980 10854 7032 10906
rect 7044 10854 7096 10906
rect 8765 10854 8817 10906
rect 8829 10854 8881 10906
rect 8893 10854 8945 10906
rect 8957 10854 9009 10906
rect 9021 10854 9073 10906
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 8392 10616 8444 10668
rect 8576 10412 8628 10464
rect 1846 10310 1898 10362
rect 1910 10310 1962 10362
rect 1974 10310 2026 10362
rect 2038 10310 2090 10362
rect 2102 10310 2154 10362
rect 3823 10310 3875 10362
rect 3887 10310 3939 10362
rect 3951 10310 4003 10362
rect 4015 10310 4067 10362
rect 4079 10310 4131 10362
rect 5800 10310 5852 10362
rect 5864 10310 5916 10362
rect 5928 10310 5980 10362
rect 5992 10310 6044 10362
rect 6056 10310 6108 10362
rect 7777 10310 7829 10362
rect 7841 10310 7893 10362
rect 7905 10310 7957 10362
rect 7969 10310 8021 10362
rect 8033 10310 8085 10362
rect 2834 9766 2886 9818
rect 2898 9766 2950 9818
rect 2962 9766 3014 9818
rect 3026 9766 3078 9818
rect 3090 9766 3142 9818
rect 4811 9766 4863 9818
rect 4875 9766 4927 9818
rect 4939 9766 4991 9818
rect 5003 9766 5055 9818
rect 5067 9766 5119 9818
rect 6788 9766 6840 9818
rect 6852 9766 6904 9818
rect 6916 9766 6968 9818
rect 6980 9766 7032 9818
rect 7044 9766 7096 9818
rect 8765 9766 8817 9818
rect 8829 9766 8881 9818
rect 8893 9766 8945 9818
rect 8957 9766 9009 9818
rect 9021 9766 9073 9818
rect 1846 9222 1898 9274
rect 1910 9222 1962 9274
rect 1974 9222 2026 9274
rect 2038 9222 2090 9274
rect 2102 9222 2154 9274
rect 3823 9222 3875 9274
rect 3887 9222 3939 9274
rect 3951 9222 4003 9274
rect 4015 9222 4067 9274
rect 4079 9222 4131 9274
rect 5800 9222 5852 9274
rect 5864 9222 5916 9274
rect 5928 9222 5980 9274
rect 5992 9222 6044 9274
rect 6056 9222 6108 9274
rect 7777 9222 7829 9274
rect 7841 9222 7893 9274
rect 7905 9222 7957 9274
rect 7969 9222 8021 9274
rect 8033 9222 8085 9274
rect 8392 8916 8444 8968
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8300 8780 8352 8832
rect 8576 8848 8628 8900
rect 2834 8678 2886 8730
rect 2898 8678 2950 8730
rect 2962 8678 3014 8730
rect 3026 8678 3078 8730
rect 3090 8678 3142 8730
rect 4811 8678 4863 8730
rect 4875 8678 4927 8730
rect 4939 8678 4991 8730
rect 5003 8678 5055 8730
rect 5067 8678 5119 8730
rect 6788 8678 6840 8730
rect 6852 8678 6904 8730
rect 6916 8678 6968 8730
rect 6980 8678 7032 8730
rect 7044 8678 7096 8730
rect 8765 8678 8817 8730
rect 8829 8678 8881 8730
rect 8893 8678 8945 8730
rect 8957 8678 9009 8730
rect 9021 8678 9073 8730
rect 1846 8134 1898 8186
rect 1910 8134 1962 8186
rect 1974 8134 2026 8186
rect 2038 8134 2090 8186
rect 2102 8134 2154 8186
rect 3823 8134 3875 8186
rect 3887 8134 3939 8186
rect 3951 8134 4003 8186
rect 4015 8134 4067 8186
rect 4079 8134 4131 8186
rect 5800 8134 5852 8186
rect 5864 8134 5916 8186
rect 5928 8134 5980 8186
rect 5992 8134 6044 8186
rect 6056 8134 6108 8186
rect 7777 8134 7829 8186
rect 7841 8134 7893 8186
rect 7905 8134 7957 8186
rect 7969 8134 8021 8186
rect 8033 8134 8085 8186
rect 2834 7590 2886 7642
rect 2898 7590 2950 7642
rect 2962 7590 3014 7642
rect 3026 7590 3078 7642
rect 3090 7590 3142 7642
rect 4811 7590 4863 7642
rect 4875 7590 4927 7642
rect 4939 7590 4991 7642
rect 5003 7590 5055 7642
rect 5067 7590 5119 7642
rect 6788 7590 6840 7642
rect 6852 7590 6904 7642
rect 6916 7590 6968 7642
rect 6980 7590 7032 7642
rect 7044 7590 7096 7642
rect 8765 7590 8817 7642
rect 8829 7590 8881 7642
rect 8893 7590 8945 7642
rect 8957 7590 9009 7642
rect 9021 7590 9073 7642
rect 1846 7046 1898 7098
rect 1910 7046 1962 7098
rect 1974 7046 2026 7098
rect 2038 7046 2090 7098
rect 2102 7046 2154 7098
rect 3823 7046 3875 7098
rect 3887 7046 3939 7098
rect 3951 7046 4003 7098
rect 4015 7046 4067 7098
rect 4079 7046 4131 7098
rect 5800 7046 5852 7098
rect 5864 7046 5916 7098
rect 5928 7046 5980 7098
rect 5992 7046 6044 7098
rect 6056 7046 6108 7098
rect 7777 7046 7829 7098
rect 7841 7046 7893 7098
rect 7905 7046 7957 7098
rect 7969 7046 8021 7098
rect 8033 7046 8085 7098
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 2834 6502 2886 6554
rect 2898 6502 2950 6554
rect 2962 6502 3014 6554
rect 3026 6502 3078 6554
rect 3090 6502 3142 6554
rect 4811 6502 4863 6554
rect 4875 6502 4927 6554
rect 4939 6502 4991 6554
rect 5003 6502 5055 6554
rect 5067 6502 5119 6554
rect 6788 6502 6840 6554
rect 6852 6502 6904 6554
rect 6916 6502 6968 6554
rect 6980 6502 7032 6554
rect 7044 6502 7096 6554
rect 8765 6502 8817 6554
rect 8829 6502 8881 6554
rect 8893 6502 8945 6554
rect 8957 6502 9009 6554
rect 9021 6502 9073 6554
rect 1846 5958 1898 6010
rect 1910 5958 1962 6010
rect 1974 5958 2026 6010
rect 2038 5958 2090 6010
rect 2102 5958 2154 6010
rect 3823 5958 3875 6010
rect 3887 5958 3939 6010
rect 3951 5958 4003 6010
rect 4015 5958 4067 6010
rect 4079 5958 4131 6010
rect 5800 5958 5852 6010
rect 5864 5958 5916 6010
rect 5928 5958 5980 6010
rect 5992 5958 6044 6010
rect 6056 5958 6108 6010
rect 7777 5958 7829 6010
rect 7841 5958 7893 6010
rect 7905 5958 7957 6010
rect 7969 5958 8021 6010
rect 8033 5958 8085 6010
rect 2834 5414 2886 5466
rect 2898 5414 2950 5466
rect 2962 5414 3014 5466
rect 3026 5414 3078 5466
rect 3090 5414 3142 5466
rect 4811 5414 4863 5466
rect 4875 5414 4927 5466
rect 4939 5414 4991 5466
rect 5003 5414 5055 5466
rect 5067 5414 5119 5466
rect 6788 5414 6840 5466
rect 6852 5414 6904 5466
rect 6916 5414 6968 5466
rect 6980 5414 7032 5466
rect 7044 5414 7096 5466
rect 8765 5414 8817 5466
rect 8829 5414 8881 5466
rect 8893 5414 8945 5466
rect 8957 5414 9009 5466
rect 9021 5414 9073 5466
rect 8392 5244 8444 5296
rect 8300 5040 8352 5092
rect 8208 4972 8260 5024
rect 1846 4870 1898 4922
rect 1910 4870 1962 4922
rect 1974 4870 2026 4922
rect 2038 4870 2090 4922
rect 2102 4870 2154 4922
rect 3823 4870 3875 4922
rect 3887 4870 3939 4922
rect 3951 4870 4003 4922
rect 4015 4870 4067 4922
rect 4079 4870 4131 4922
rect 5800 4870 5852 4922
rect 5864 4870 5916 4922
rect 5928 4870 5980 4922
rect 5992 4870 6044 4922
rect 6056 4870 6108 4922
rect 7777 4870 7829 4922
rect 7841 4870 7893 4922
rect 7905 4870 7957 4922
rect 7969 4870 8021 4922
rect 8033 4870 8085 4922
rect 2834 4326 2886 4378
rect 2898 4326 2950 4378
rect 2962 4326 3014 4378
rect 3026 4326 3078 4378
rect 3090 4326 3142 4378
rect 4811 4326 4863 4378
rect 4875 4326 4927 4378
rect 4939 4326 4991 4378
rect 5003 4326 5055 4378
rect 5067 4326 5119 4378
rect 6788 4326 6840 4378
rect 6852 4326 6904 4378
rect 6916 4326 6968 4378
rect 6980 4326 7032 4378
rect 7044 4326 7096 4378
rect 8765 4326 8817 4378
rect 8829 4326 8881 4378
rect 8893 4326 8945 4378
rect 8957 4326 9009 4378
rect 9021 4326 9073 4378
rect 1846 3782 1898 3834
rect 1910 3782 1962 3834
rect 1974 3782 2026 3834
rect 2038 3782 2090 3834
rect 2102 3782 2154 3834
rect 3823 3782 3875 3834
rect 3887 3782 3939 3834
rect 3951 3782 4003 3834
rect 4015 3782 4067 3834
rect 4079 3782 4131 3834
rect 5800 3782 5852 3834
rect 5864 3782 5916 3834
rect 5928 3782 5980 3834
rect 5992 3782 6044 3834
rect 6056 3782 6108 3834
rect 7777 3782 7829 3834
rect 7841 3782 7893 3834
rect 7905 3782 7957 3834
rect 7969 3782 8021 3834
rect 8033 3782 8085 3834
rect 2834 3238 2886 3290
rect 2898 3238 2950 3290
rect 2962 3238 3014 3290
rect 3026 3238 3078 3290
rect 3090 3238 3142 3290
rect 4811 3238 4863 3290
rect 4875 3238 4927 3290
rect 4939 3238 4991 3290
rect 5003 3238 5055 3290
rect 5067 3238 5119 3290
rect 6788 3238 6840 3290
rect 6852 3238 6904 3290
rect 6916 3238 6968 3290
rect 6980 3238 7032 3290
rect 7044 3238 7096 3290
rect 8765 3238 8817 3290
rect 8829 3238 8881 3290
rect 8893 3238 8945 3290
rect 8957 3238 9009 3290
rect 9021 3238 9073 3290
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 8300 3000 8352 3052
rect 8116 2907 8168 2916
rect 8116 2873 8125 2907
rect 8125 2873 8159 2907
rect 8159 2873 8168 2907
rect 8116 2864 8168 2873
rect 8300 2864 8352 2916
rect 8392 2796 8444 2848
rect 1846 2694 1898 2746
rect 1910 2694 1962 2746
rect 1974 2694 2026 2746
rect 2038 2694 2090 2746
rect 2102 2694 2154 2746
rect 3823 2694 3875 2746
rect 3887 2694 3939 2746
rect 3951 2694 4003 2746
rect 4015 2694 4067 2746
rect 4079 2694 4131 2746
rect 5800 2694 5852 2746
rect 5864 2694 5916 2746
rect 5928 2694 5980 2746
rect 5992 2694 6044 2746
rect 6056 2694 6108 2746
rect 7777 2694 7829 2746
rect 7841 2694 7893 2746
rect 7905 2694 7957 2746
rect 7969 2694 8021 2746
rect 8033 2694 8085 2746
rect 2834 2150 2886 2202
rect 2898 2150 2950 2202
rect 2962 2150 3014 2202
rect 3026 2150 3078 2202
rect 3090 2150 3142 2202
rect 4811 2150 4863 2202
rect 4875 2150 4927 2202
rect 4939 2150 4991 2202
rect 5003 2150 5055 2202
rect 5067 2150 5119 2202
rect 6788 2150 6840 2202
rect 6852 2150 6904 2202
rect 6916 2150 6968 2202
rect 6980 2150 7032 2202
rect 7044 2150 7096 2202
rect 8765 2150 8817 2202
rect 8829 2150 8881 2202
rect 8893 2150 8945 2202
rect 8957 2150 9009 2202
rect 9021 2150 9073 2202
rect 8116 1955 8168 1964
rect 8116 1921 8125 1955
rect 8125 1921 8159 1955
rect 8159 1921 8168 1955
rect 8116 1912 8168 1921
rect 8300 1955 8352 1964
rect 8300 1921 8309 1955
rect 8309 1921 8343 1955
rect 8343 1921 8352 1955
rect 8300 1912 8352 1921
rect 9312 1844 9364 1896
rect 1846 1606 1898 1658
rect 1910 1606 1962 1658
rect 1974 1606 2026 1658
rect 2038 1606 2090 1658
rect 2102 1606 2154 1658
rect 3823 1606 3875 1658
rect 3887 1606 3939 1658
rect 3951 1606 4003 1658
rect 4015 1606 4067 1658
rect 4079 1606 4131 1658
rect 5800 1606 5852 1658
rect 5864 1606 5916 1658
rect 5928 1606 5980 1658
rect 5992 1606 6044 1658
rect 6056 1606 6108 1658
rect 7777 1606 7829 1658
rect 7841 1606 7893 1658
rect 7905 1606 7957 1658
rect 7969 1606 8021 1658
rect 8033 1606 8085 1658
rect 8116 1504 8168 1556
rect 8300 1436 8352 1488
rect 7472 1300 7524 1352
rect 2504 1232 2556 1284
rect 2834 1062 2886 1114
rect 2898 1062 2950 1114
rect 2962 1062 3014 1114
rect 3026 1062 3078 1114
rect 3090 1062 3142 1114
rect 4811 1062 4863 1114
rect 4875 1062 4927 1114
rect 4939 1062 4991 1114
rect 5003 1062 5055 1114
rect 5067 1062 5119 1114
rect 6788 1062 6840 1114
rect 6852 1062 6904 1114
rect 6916 1062 6968 1114
rect 6980 1062 7032 1114
rect 7044 1062 7096 1114
rect 8765 1062 8817 1114
rect 8829 1062 8881 1114
rect 8893 1062 8945 1114
rect 8957 1062 9009 1114
rect 9021 1062 9073 1114
<< metal2 >>
rect 1846 14716 2154 14725
rect 1846 14714 1852 14716
rect 1908 14714 1932 14716
rect 1988 14714 2012 14716
rect 2068 14714 2092 14716
rect 2148 14714 2154 14716
rect 1908 14662 1910 14714
rect 2090 14662 2092 14714
rect 1846 14660 1852 14662
rect 1908 14660 1932 14662
rect 1988 14660 2012 14662
rect 2068 14660 2092 14662
rect 2148 14660 2154 14662
rect 1846 14651 2154 14660
rect 3823 14716 4131 14725
rect 3823 14714 3829 14716
rect 3885 14714 3909 14716
rect 3965 14714 3989 14716
rect 4045 14714 4069 14716
rect 4125 14714 4131 14716
rect 3885 14662 3887 14714
rect 4067 14662 4069 14714
rect 3823 14660 3829 14662
rect 3885 14660 3909 14662
rect 3965 14660 3989 14662
rect 4045 14660 4069 14662
rect 4125 14660 4131 14662
rect 3823 14651 4131 14660
rect 5800 14716 6108 14725
rect 5800 14714 5806 14716
rect 5862 14714 5886 14716
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6108 14716
rect 5862 14662 5864 14714
rect 6044 14662 6046 14714
rect 5800 14660 5806 14662
rect 5862 14660 5886 14662
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6108 14662
rect 5800 14651 6108 14660
rect 7777 14716 8085 14725
rect 7777 14714 7783 14716
rect 7839 14714 7863 14716
rect 7919 14714 7943 14716
rect 7999 14714 8023 14716
rect 8079 14714 8085 14716
rect 7839 14662 7841 14714
rect 8021 14662 8023 14714
rect 7777 14660 7783 14662
rect 7839 14660 7863 14662
rect 7919 14660 7943 14662
rect 7999 14660 8023 14662
rect 8079 14660 8085 14662
rect 7777 14651 8085 14660
rect 8114 14512 8170 14521
rect 8114 14447 8170 14456
rect 2834 14172 3142 14181
rect 2834 14170 2840 14172
rect 2896 14170 2920 14172
rect 2976 14170 3000 14172
rect 3056 14170 3080 14172
rect 3136 14170 3142 14172
rect 2896 14118 2898 14170
rect 3078 14118 3080 14170
rect 2834 14116 2840 14118
rect 2896 14116 2920 14118
rect 2976 14116 3000 14118
rect 3056 14116 3080 14118
rect 3136 14116 3142 14118
rect 2834 14107 3142 14116
rect 4811 14172 5119 14181
rect 4811 14170 4817 14172
rect 4873 14170 4897 14172
rect 4953 14170 4977 14172
rect 5033 14170 5057 14172
rect 5113 14170 5119 14172
rect 4873 14118 4875 14170
rect 5055 14118 5057 14170
rect 4811 14116 4817 14118
rect 4873 14116 4897 14118
rect 4953 14116 4977 14118
rect 5033 14116 5057 14118
rect 5113 14116 5119 14118
rect 4811 14107 5119 14116
rect 6788 14172 7096 14181
rect 6788 14170 6794 14172
rect 6850 14170 6874 14172
rect 6930 14170 6954 14172
rect 7010 14170 7034 14172
rect 7090 14170 7096 14172
rect 6850 14118 6852 14170
rect 7032 14118 7034 14170
rect 6788 14116 6794 14118
rect 6850 14116 6874 14118
rect 6930 14116 6954 14118
rect 7010 14116 7034 14118
rect 7090 14116 7096 14118
rect 6788 14107 7096 14116
rect 1846 13628 2154 13637
rect 1846 13626 1852 13628
rect 1908 13626 1932 13628
rect 1988 13626 2012 13628
rect 2068 13626 2092 13628
rect 2148 13626 2154 13628
rect 1908 13574 1910 13626
rect 2090 13574 2092 13626
rect 1846 13572 1852 13574
rect 1908 13572 1932 13574
rect 1988 13572 2012 13574
rect 2068 13572 2092 13574
rect 2148 13572 2154 13574
rect 1846 13563 2154 13572
rect 3823 13628 4131 13637
rect 3823 13626 3829 13628
rect 3885 13626 3909 13628
rect 3965 13626 3989 13628
rect 4045 13626 4069 13628
rect 4125 13626 4131 13628
rect 3885 13574 3887 13626
rect 4067 13574 4069 13626
rect 3823 13572 3829 13574
rect 3885 13572 3909 13574
rect 3965 13572 3989 13574
rect 4045 13572 4069 13574
rect 4125 13572 4131 13574
rect 3823 13563 4131 13572
rect 5800 13628 6108 13637
rect 5800 13626 5806 13628
rect 5862 13626 5886 13628
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6108 13628
rect 5862 13574 5864 13626
rect 6044 13574 6046 13626
rect 5800 13572 5806 13574
rect 5862 13572 5886 13574
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6108 13574
rect 5800 13563 6108 13572
rect 7777 13628 8085 13637
rect 7777 13626 7783 13628
rect 7839 13626 7863 13628
rect 7919 13626 7943 13628
rect 7999 13626 8023 13628
rect 8079 13626 8085 13628
rect 7839 13574 7841 13626
rect 8021 13574 8023 13626
rect 7777 13572 7783 13574
rect 7839 13572 7863 13574
rect 7919 13572 7943 13574
rect 7999 13572 8023 13574
rect 8079 13572 8085 13574
rect 7777 13563 8085 13572
rect 2834 13084 3142 13093
rect 2834 13082 2840 13084
rect 2896 13082 2920 13084
rect 2976 13082 3000 13084
rect 3056 13082 3080 13084
rect 3136 13082 3142 13084
rect 2896 13030 2898 13082
rect 3078 13030 3080 13082
rect 2834 13028 2840 13030
rect 2896 13028 2920 13030
rect 2976 13028 3000 13030
rect 3056 13028 3080 13030
rect 3136 13028 3142 13030
rect 2834 13019 3142 13028
rect 4811 13084 5119 13093
rect 4811 13082 4817 13084
rect 4873 13082 4897 13084
rect 4953 13082 4977 13084
rect 5033 13082 5057 13084
rect 5113 13082 5119 13084
rect 4873 13030 4875 13082
rect 5055 13030 5057 13082
rect 4811 13028 4817 13030
rect 4873 13028 4897 13030
rect 4953 13028 4977 13030
rect 5033 13028 5057 13030
rect 5113 13028 5119 13030
rect 4811 13019 5119 13028
rect 6788 13084 7096 13093
rect 6788 13082 6794 13084
rect 6850 13082 6874 13084
rect 6930 13082 6954 13084
rect 7010 13082 7034 13084
rect 7090 13082 7096 13084
rect 6850 13030 6852 13082
rect 7032 13030 7034 13082
rect 6788 13028 6794 13030
rect 6850 13028 6874 13030
rect 6930 13028 6954 13030
rect 7010 13028 7034 13030
rect 7090 13028 7096 13030
rect 6788 13019 7096 13028
rect 1846 12540 2154 12549
rect 1846 12538 1852 12540
rect 1908 12538 1932 12540
rect 1988 12538 2012 12540
rect 2068 12538 2092 12540
rect 2148 12538 2154 12540
rect 1908 12486 1910 12538
rect 2090 12486 2092 12538
rect 1846 12484 1852 12486
rect 1908 12484 1932 12486
rect 1988 12484 2012 12486
rect 2068 12484 2092 12486
rect 2148 12484 2154 12486
rect 1846 12475 2154 12484
rect 3823 12540 4131 12549
rect 3823 12538 3829 12540
rect 3885 12538 3909 12540
rect 3965 12538 3989 12540
rect 4045 12538 4069 12540
rect 4125 12538 4131 12540
rect 3885 12486 3887 12538
rect 4067 12486 4069 12538
rect 3823 12484 3829 12486
rect 3885 12484 3909 12486
rect 3965 12484 3989 12486
rect 4045 12484 4069 12486
rect 4125 12484 4131 12486
rect 3823 12475 4131 12484
rect 5800 12540 6108 12549
rect 5800 12538 5806 12540
rect 5862 12538 5886 12540
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6108 12540
rect 5862 12486 5864 12538
rect 6044 12486 6046 12538
rect 5800 12484 5806 12486
rect 5862 12484 5886 12486
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6108 12486
rect 5800 12475 6108 12484
rect 7777 12540 8085 12549
rect 7777 12538 7783 12540
rect 7839 12538 7863 12540
rect 7919 12538 7943 12540
rect 7999 12538 8023 12540
rect 8079 12538 8085 12540
rect 7839 12486 7841 12538
rect 8021 12486 8023 12538
rect 7777 12484 7783 12486
rect 7839 12484 7863 12486
rect 7919 12484 7943 12486
rect 7999 12484 8023 12486
rect 8079 12484 8085 12486
rect 7777 12475 8085 12484
rect 2834 11996 3142 12005
rect 2834 11994 2840 11996
rect 2896 11994 2920 11996
rect 2976 11994 3000 11996
rect 3056 11994 3080 11996
rect 3136 11994 3142 11996
rect 2896 11942 2898 11994
rect 3078 11942 3080 11994
rect 2834 11940 2840 11942
rect 2896 11940 2920 11942
rect 2976 11940 3000 11942
rect 3056 11940 3080 11942
rect 3136 11940 3142 11942
rect 2834 11931 3142 11940
rect 4811 11996 5119 12005
rect 4811 11994 4817 11996
rect 4873 11994 4897 11996
rect 4953 11994 4977 11996
rect 5033 11994 5057 11996
rect 5113 11994 5119 11996
rect 4873 11942 4875 11994
rect 5055 11942 5057 11994
rect 4811 11940 4817 11942
rect 4873 11940 4897 11942
rect 4953 11940 4977 11942
rect 5033 11940 5057 11942
rect 5113 11940 5119 11942
rect 4811 11931 5119 11940
rect 6788 11996 7096 12005
rect 6788 11994 6794 11996
rect 6850 11994 6874 11996
rect 6930 11994 6954 11996
rect 7010 11994 7034 11996
rect 7090 11994 7096 11996
rect 6850 11942 6852 11994
rect 7032 11942 7034 11994
rect 6788 11940 6794 11942
rect 6850 11940 6874 11942
rect 6930 11940 6954 11942
rect 7010 11940 7034 11942
rect 7090 11940 7096 11942
rect 6788 11931 7096 11940
rect 8128 11762 8156 14447
rect 8765 14172 9073 14181
rect 8765 14170 8771 14172
rect 8827 14170 8851 14172
rect 8907 14170 8931 14172
rect 8987 14170 9011 14172
rect 9067 14170 9073 14172
rect 8827 14118 8829 14170
rect 9009 14118 9011 14170
rect 8765 14116 8771 14118
rect 8827 14116 8851 14118
rect 8907 14116 8931 14118
rect 8987 14116 9011 14118
rect 9067 14116 9073 14118
rect 8765 14107 9073 14116
rect 8765 13084 9073 13093
rect 8765 13082 8771 13084
rect 8827 13082 8851 13084
rect 8907 13082 8931 13084
rect 8987 13082 9011 13084
rect 9067 13082 9073 13084
rect 8827 13030 8829 13082
rect 9009 13030 9011 13082
rect 8765 13028 8771 13030
rect 8827 13028 8851 13030
rect 8907 13028 8931 13030
rect 8987 13028 9011 13030
rect 9067 13028 9073 13030
rect 8765 13019 9073 13028
rect 8206 12608 8262 12617
rect 8206 12543 8262 12552
rect 8220 12442 8248 12543
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 1846 11452 2154 11461
rect 1846 11450 1852 11452
rect 1908 11450 1932 11452
rect 1988 11450 2012 11452
rect 2068 11450 2092 11452
rect 2148 11450 2154 11452
rect 1908 11398 1910 11450
rect 2090 11398 2092 11450
rect 1846 11396 1852 11398
rect 1908 11396 1932 11398
rect 1988 11396 2012 11398
rect 2068 11396 2092 11398
rect 2148 11396 2154 11398
rect 1846 11387 2154 11396
rect 3823 11452 4131 11461
rect 3823 11450 3829 11452
rect 3885 11450 3909 11452
rect 3965 11450 3989 11452
rect 4045 11450 4069 11452
rect 4125 11450 4131 11452
rect 3885 11398 3887 11450
rect 4067 11398 4069 11450
rect 3823 11396 3829 11398
rect 3885 11396 3909 11398
rect 3965 11396 3989 11398
rect 4045 11396 4069 11398
rect 4125 11396 4131 11398
rect 3823 11387 4131 11396
rect 5800 11452 6108 11461
rect 5800 11450 5806 11452
rect 5862 11450 5886 11452
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6108 11452
rect 5862 11398 5864 11450
rect 6044 11398 6046 11450
rect 5800 11396 5806 11398
rect 5862 11396 5886 11398
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6108 11398
rect 5800 11387 6108 11396
rect 7777 11452 8085 11461
rect 7777 11450 7783 11452
rect 7839 11450 7863 11452
rect 7919 11450 7943 11452
rect 7999 11450 8023 11452
rect 8079 11450 8085 11452
rect 7839 11398 7841 11450
rect 8021 11398 8023 11450
rect 7777 11396 7783 11398
rect 7839 11396 7863 11398
rect 7919 11396 7943 11398
rect 7999 11396 8023 11398
rect 8079 11396 8085 11398
rect 7777 11387 8085 11396
rect 8404 11354 8432 11630
rect 8496 11354 8524 12174
rect 8765 11996 9073 12005
rect 8765 11994 8771 11996
rect 8827 11994 8851 11996
rect 8907 11994 8931 11996
rect 8987 11994 9011 11996
rect 9067 11994 9073 11996
rect 8827 11942 8829 11994
rect 9009 11942 9011 11994
rect 8765 11940 8771 11942
rect 8827 11940 8851 11942
rect 8907 11940 8931 11942
rect 8987 11940 9011 11942
rect 9067 11940 9073 11942
rect 8765 11931 9073 11940
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 2834 10908 3142 10917
rect 2834 10906 2840 10908
rect 2896 10906 2920 10908
rect 2976 10906 3000 10908
rect 3056 10906 3080 10908
rect 3136 10906 3142 10908
rect 2896 10854 2898 10906
rect 3078 10854 3080 10906
rect 2834 10852 2840 10854
rect 2896 10852 2920 10854
rect 2976 10852 3000 10854
rect 3056 10852 3080 10854
rect 3136 10852 3142 10854
rect 2834 10843 3142 10852
rect 4811 10908 5119 10917
rect 4811 10906 4817 10908
rect 4873 10906 4897 10908
rect 4953 10906 4977 10908
rect 5033 10906 5057 10908
rect 5113 10906 5119 10908
rect 4873 10854 4875 10906
rect 5055 10854 5057 10906
rect 4811 10852 4817 10854
rect 4873 10852 4897 10854
rect 4953 10852 4977 10854
rect 5033 10852 5057 10854
rect 5113 10852 5119 10854
rect 4811 10843 5119 10852
rect 6788 10908 7096 10917
rect 6788 10906 6794 10908
rect 6850 10906 6874 10908
rect 6930 10906 6954 10908
rect 7010 10906 7034 10908
rect 7090 10906 7096 10908
rect 6850 10854 6852 10906
rect 7032 10854 7034 10906
rect 6788 10852 6794 10854
rect 6850 10852 6874 10854
rect 6930 10852 6954 10854
rect 7010 10852 7034 10854
rect 7090 10852 7096 10854
rect 6788 10843 7096 10852
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7760 10713 7788 10746
rect 7746 10704 7802 10713
rect 8404 10674 8432 11290
rect 8588 11150 8616 11698
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 7746 10639 7802 10648
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 1846 10364 2154 10373
rect 1846 10362 1852 10364
rect 1908 10362 1932 10364
rect 1988 10362 2012 10364
rect 2068 10362 2092 10364
rect 2148 10362 2154 10364
rect 1908 10310 1910 10362
rect 2090 10310 2092 10362
rect 1846 10308 1852 10310
rect 1908 10308 1932 10310
rect 1988 10308 2012 10310
rect 2068 10308 2092 10310
rect 2148 10308 2154 10310
rect 1846 10299 2154 10308
rect 3823 10364 4131 10373
rect 3823 10362 3829 10364
rect 3885 10362 3909 10364
rect 3965 10362 3989 10364
rect 4045 10362 4069 10364
rect 4125 10362 4131 10364
rect 3885 10310 3887 10362
rect 4067 10310 4069 10362
rect 3823 10308 3829 10310
rect 3885 10308 3909 10310
rect 3965 10308 3989 10310
rect 4045 10308 4069 10310
rect 4125 10308 4131 10310
rect 3823 10299 4131 10308
rect 5800 10364 6108 10373
rect 5800 10362 5806 10364
rect 5862 10362 5886 10364
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6108 10364
rect 5862 10310 5864 10362
rect 6044 10310 6046 10362
rect 5800 10308 5806 10310
rect 5862 10308 5886 10310
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6108 10310
rect 5800 10299 6108 10308
rect 7777 10364 8085 10373
rect 7777 10362 7783 10364
rect 7839 10362 7863 10364
rect 7919 10362 7943 10364
rect 7999 10362 8023 10364
rect 8079 10362 8085 10364
rect 7839 10310 7841 10362
rect 8021 10310 8023 10362
rect 7777 10308 7783 10310
rect 7839 10308 7863 10310
rect 7919 10308 7943 10310
rect 7999 10308 8023 10310
rect 8079 10308 8085 10310
rect 7777 10299 8085 10308
rect 2834 9820 3142 9829
rect 2834 9818 2840 9820
rect 2896 9818 2920 9820
rect 2976 9818 3000 9820
rect 3056 9818 3080 9820
rect 3136 9818 3142 9820
rect 2896 9766 2898 9818
rect 3078 9766 3080 9818
rect 2834 9764 2840 9766
rect 2896 9764 2920 9766
rect 2976 9764 3000 9766
rect 3056 9764 3080 9766
rect 3136 9764 3142 9766
rect 2834 9755 3142 9764
rect 4811 9820 5119 9829
rect 4811 9818 4817 9820
rect 4873 9818 4897 9820
rect 4953 9818 4977 9820
rect 5033 9818 5057 9820
rect 5113 9818 5119 9820
rect 4873 9766 4875 9818
rect 5055 9766 5057 9818
rect 4811 9764 4817 9766
rect 4873 9764 4897 9766
rect 4953 9764 4977 9766
rect 5033 9764 5057 9766
rect 5113 9764 5119 9766
rect 4811 9755 5119 9764
rect 6788 9820 7096 9829
rect 6788 9818 6794 9820
rect 6850 9818 6874 9820
rect 6930 9818 6954 9820
rect 7010 9818 7034 9820
rect 7090 9818 7096 9820
rect 6850 9766 6852 9818
rect 7032 9766 7034 9818
rect 6788 9764 6794 9766
rect 6850 9764 6874 9766
rect 6930 9764 6954 9766
rect 7010 9764 7034 9766
rect 7090 9764 7096 9766
rect 6788 9755 7096 9764
rect 1846 9276 2154 9285
rect 1846 9274 1852 9276
rect 1908 9274 1932 9276
rect 1988 9274 2012 9276
rect 2068 9274 2092 9276
rect 2148 9274 2154 9276
rect 1908 9222 1910 9274
rect 2090 9222 2092 9274
rect 1846 9220 1852 9222
rect 1908 9220 1932 9222
rect 1988 9220 2012 9222
rect 2068 9220 2092 9222
rect 2148 9220 2154 9222
rect 1846 9211 2154 9220
rect 3823 9276 4131 9285
rect 3823 9274 3829 9276
rect 3885 9274 3909 9276
rect 3965 9274 3989 9276
rect 4045 9274 4069 9276
rect 4125 9274 4131 9276
rect 3885 9222 3887 9274
rect 4067 9222 4069 9274
rect 3823 9220 3829 9222
rect 3885 9220 3909 9222
rect 3965 9220 3989 9222
rect 4045 9220 4069 9222
rect 4125 9220 4131 9222
rect 3823 9211 4131 9220
rect 5800 9276 6108 9285
rect 5800 9274 5806 9276
rect 5862 9274 5886 9276
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6108 9276
rect 5862 9222 5864 9274
rect 6044 9222 6046 9274
rect 5800 9220 5806 9222
rect 5862 9220 5886 9222
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6108 9222
rect 5800 9211 6108 9220
rect 7777 9276 8085 9285
rect 7777 9274 7783 9276
rect 7839 9274 7863 9276
rect 7919 9274 7943 9276
rect 7999 9274 8023 9276
rect 8079 9274 8085 9276
rect 7839 9222 7841 9274
rect 8021 9222 8023 9274
rect 7777 9220 7783 9222
rect 7839 9220 7863 9222
rect 7919 9220 7943 9222
rect 7999 9220 8023 9222
rect 8079 9220 8085 9222
rect 7777 9211 8085 9220
rect 8404 8974 8432 10610
rect 8588 10470 8616 11086
rect 8765 10908 9073 10917
rect 8765 10906 8771 10908
rect 8827 10906 8851 10908
rect 8907 10906 8931 10908
rect 8987 10906 9011 10908
rect 9067 10906 9073 10908
rect 8827 10854 8829 10906
rect 9009 10854 9011 10906
rect 8765 10852 8771 10854
rect 8827 10852 8851 10854
rect 8907 10852 8931 10854
rect 8987 10852 9011 10854
rect 9067 10852 9073 10854
rect 8765 10843 9073 10852
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8392 8968 8444 8974
rect 7838 8936 7894 8945
rect 8392 8910 8444 8916
rect 7838 8871 7894 8880
rect 7852 8838 7880 8871
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 2834 8732 3142 8741
rect 2834 8730 2840 8732
rect 2896 8730 2920 8732
rect 2976 8730 3000 8732
rect 3056 8730 3080 8732
rect 3136 8730 3142 8732
rect 2896 8678 2898 8730
rect 3078 8678 3080 8730
rect 2834 8676 2840 8678
rect 2896 8676 2920 8678
rect 2976 8676 3000 8678
rect 3056 8676 3080 8678
rect 3136 8676 3142 8678
rect 2834 8667 3142 8676
rect 4811 8732 5119 8741
rect 4811 8730 4817 8732
rect 4873 8730 4897 8732
rect 4953 8730 4977 8732
rect 5033 8730 5057 8732
rect 5113 8730 5119 8732
rect 4873 8678 4875 8730
rect 5055 8678 5057 8730
rect 4811 8676 4817 8678
rect 4873 8676 4897 8678
rect 4953 8676 4977 8678
rect 5033 8676 5057 8678
rect 5113 8676 5119 8678
rect 4811 8667 5119 8676
rect 6788 8732 7096 8741
rect 6788 8730 6794 8732
rect 6850 8730 6874 8732
rect 6930 8730 6954 8732
rect 7010 8730 7034 8732
rect 7090 8730 7096 8732
rect 6850 8678 6852 8730
rect 7032 8678 7034 8730
rect 6788 8676 6794 8678
rect 6850 8676 6874 8678
rect 6930 8676 6954 8678
rect 7010 8676 7034 8678
rect 7090 8676 7096 8678
rect 6788 8667 7096 8676
rect 1846 8188 2154 8197
rect 1846 8186 1852 8188
rect 1908 8186 1932 8188
rect 1988 8186 2012 8188
rect 2068 8186 2092 8188
rect 2148 8186 2154 8188
rect 1908 8134 1910 8186
rect 2090 8134 2092 8186
rect 1846 8132 1852 8134
rect 1908 8132 1932 8134
rect 1988 8132 2012 8134
rect 2068 8132 2092 8134
rect 2148 8132 2154 8134
rect 1846 8123 2154 8132
rect 3823 8188 4131 8197
rect 3823 8186 3829 8188
rect 3885 8186 3909 8188
rect 3965 8186 3989 8188
rect 4045 8186 4069 8188
rect 4125 8186 4131 8188
rect 3885 8134 3887 8186
rect 4067 8134 4069 8186
rect 3823 8132 3829 8134
rect 3885 8132 3909 8134
rect 3965 8132 3989 8134
rect 4045 8132 4069 8134
rect 4125 8132 4131 8134
rect 3823 8123 4131 8132
rect 5800 8188 6108 8197
rect 5800 8186 5806 8188
rect 5862 8186 5886 8188
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6108 8188
rect 5862 8134 5864 8186
rect 6044 8134 6046 8186
rect 5800 8132 5806 8134
rect 5862 8132 5886 8134
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6108 8134
rect 5800 8123 6108 8132
rect 7777 8188 8085 8197
rect 7777 8186 7783 8188
rect 7839 8186 7863 8188
rect 7919 8186 7943 8188
rect 7999 8186 8023 8188
rect 8079 8186 8085 8188
rect 7839 8134 7841 8186
rect 8021 8134 8023 8186
rect 7777 8132 7783 8134
rect 7839 8132 7863 8134
rect 7919 8132 7943 8134
rect 7999 8132 8023 8134
rect 8079 8132 8085 8134
rect 7777 8123 8085 8132
rect 2834 7644 3142 7653
rect 2834 7642 2840 7644
rect 2896 7642 2920 7644
rect 2976 7642 3000 7644
rect 3056 7642 3080 7644
rect 3136 7642 3142 7644
rect 2896 7590 2898 7642
rect 3078 7590 3080 7642
rect 2834 7588 2840 7590
rect 2896 7588 2920 7590
rect 2976 7588 3000 7590
rect 3056 7588 3080 7590
rect 3136 7588 3142 7590
rect 2834 7579 3142 7588
rect 4811 7644 5119 7653
rect 4811 7642 4817 7644
rect 4873 7642 4897 7644
rect 4953 7642 4977 7644
rect 5033 7642 5057 7644
rect 5113 7642 5119 7644
rect 4873 7590 4875 7642
rect 5055 7590 5057 7642
rect 4811 7588 4817 7590
rect 4873 7588 4897 7590
rect 4953 7588 4977 7590
rect 5033 7588 5057 7590
rect 5113 7588 5119 7590
rect 4811 7579 5119 7588
rect 6788 7644 7096 7653
rect 6788 7642 6794 7644
rect 6850 7642 6874 7644
rect 6930 7642 6954 7644
rect 7010 7642 7034 7644
rect 7090 7642 7096 7644
rect 6850 7590 6852 7642
rect 7032 7590 7034 7642
rect 6788 7588 6794 7590
rect 6850 7588 6874 7590
rect 6930 7588 6954 7590
rect 7010 7588 7034 7590
rect 7090 7588 7096 7590
rect 6788 7579 7096 7588
rect 1846 7100 2154 7109
rect 1846 7098 1852 7100
rect 1908 7098 1932 7100
rect 1988 7098 2012 7100
rect 2068 7098 2092 7100
rect 2148 7098 2154 7100
rect 1908 7046 1910 7098
rect 2090 7046 2092 7098
rect 1846 7044 1852 7046
rect 1908 7044 1932 7046
rect 1988 7044 2012 7046
rect 2068 7044 2092 7046
rect 2148 7044 2154 7046
rect 1846 7035 2154 7044
rect 3823 7100 4131 7109
rect 3823 7098 3829 7100
rect 3885 7098 3909 7100
rect 3965 7098 3989 7100
rect 4045 7098 4069 7100
rect 4125 7098 4131 7100
rect 3885 7046 3887 7098
rect 4067 7046 4069 7098
rect 3823 7044 3829 7046
rect 3885 7044 3909 7046
rect 3965 7044 3989 7046
rect 4045 7044 4069 7046
rect 4125 7044 4131 7046
rect 3823 7035 4131 7044
rect 5800 7100 6108 7109
rect 5800 7098 5806 7100
rect 5862 7098 5886 7100
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6108 7100
rect 5862 7046 5864 7098
rect 6044 7046 6046 7098
rect 5800 7044 5806 7046
rect 5862 7044 5886 7046
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6108 7046
rect 5800 7035 6108 7044
rect 7777 7100 8085 7109
rect 7777 7098 7783 7100
rect 7839 7098 7863 7100
rect 7919 7098 7943 7100
rect 7999 7098 8023 7100
rect 8079 7098 8085 7100
rect 7839 7046 7841 7098
rect 8021 7046 8023 7098
rect 7777 7044 7783 7046
rect 7839 7044 7863 7046
rect 7919 7044 7943 7046
rect 7999 7044 8023 7046
rect 8079 7044 8085 7046
rect 7777 7035 8085 7044
rect 7838 6896 7894 6905
rect 7838 6831 7894 6840
rect 7852 6662 7880 6831
rect 8312 6798 8340 8774
rect 8404 6798 8432 8910
rect 8588 8906 8616 10406
rect 8765 9820 9073 9829
rect 8765 9818 8771 9820
rect 8827 9818 8851 9820
rect 8907 9818 8931 9820
rect 8987 9818 9011 9820
rect 9067 9818 9073 9820
rect 8827 9766 8829 9818
rect 9009 9766 9011 9818
rect 8765 9764 8771 9766
rect 8827 9764 8851 9766
rect 8907 9764 8931 9766
rect 8987 9764 9011 9766
rect 9067 9764 9073 9766
rect 8765 9755 9073 9764
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8765 8732 9073 8741
rect 8765 8730 8771 8732
rect 8827 8730 8851 8732
rect 8907 8730 8931 8732
rect 8987 8730 9011 8732
rect 9067 8730 9073 8732
rect 8827 8678 8829 8730
rect 9009 8678 9011 8730
rect 8765 8676 8771 8678
rect 8827 8676 8851 8678
rect 8907 8676 8931 8678
rect 8987 8676 9011 8678
rect 9067 8676 9073 8678
rect 8765 8667 9073 8676
rect 8765 7644 9073 7653
rect 8765 7642 8771 7644
rect 8827 7642 8851 7644
rect 8907 7642 8931 7644
rect 8987 7642 9011 7644
rect 9067 7642 9073 7644
rect 8827 7590 8829 7642
rect 9009 7590 9011 7642
rect 8765 7588 8771 7590
rect 8827 7588 8851 7590
rect 8907 7588 8931 7590
rect 8987 7588 9011 7590
rect 9067 7588 9073 7590
rect 8765 7579 9073 7588
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 2834 6556 3142 6565
rect 2834 6554 2840 6556
rect 2896 6554 2920 6556
rect 2976 6554 3000 6556
rect 3056 6554 3080 6556
rect 3136 6554 3142 6556
rect 2896 6502 2898 6554
rect 3078 6502 3080 6554
rect 2834 6500 2840 6502
rect 2896 6500 2920 6502
rect 2976 6500 3000 6502
rect 3056 6500 3080 6502
rect 3136 6500 3142 6502
rect 2834 6491 3142 6500
rect 4811 6556 5119 6565
rect 4811 6554 4817 6556
rect 4873 6554 4897 6556
rect 4953 6554 4977 6556
rect 5033 6554 5057 6556
rect 5113 6554 5119 6556
rect 4873 6502 4875 6554
rect 5055 6502 5057 6554
rect 4811 6500 4817 6502
rect 4873 6500 4897 6502
rect 4953 6500 4977 6502
rect 5033 6500 5057 6502
rect 5113 6500 5119 6502
rect 4811 6491 5119 6500
rect 6788 6556 7096 6565
rect 6788 6554 6794 6556
rect 6850 6554 6874 6556
rect 6930 6554 6954 6556
rect 7010 6554 7034 6556
rect 7090 6554 7096 6556
rect 6850 6502 6852 6554
rect 7032 6502 7034 6554
rect 6788 6500 6794 6502
rect 6850 6500 6874 6502
rect 6930 6500 6954 6502
rect 7010 6500 7034 6502
rect 7090 6500 7096 6502
rect 6788 6491 7096 6500
rect 1846 6012 2154 6021
rect 1846 6010 1852 6012
rect 1908 6010 1932 6012
rect 1988 6010 2012 6012
rect 2068 6010 2092 6012
rect 2148 6010 2154 6012
rect 1908 5958 1910 6010
rect 2090 5958 2092 6010
rect 1846 5956 1852 5958
rect 1908 5956 1932 5958
rect 1988 5956 2012 5958
rect 2068 5956 2092 5958
rect 2148 5956 2154 5958
rect 1846 5947 2154 5956
rect 3823 6012 4131 6021
rect 3823 6010 3829 6012
rect 3885 6010 3909 6012
rect 3965 6010 3989 6012
rect 4045 6010 4069 6012
rect 4125 6010 4131 6012
rect 3885 5958 3887 6010
rect 4067 5958 4069 6010
rect 3823 5956 3829 5958
rect 3885 5956 3909 5958
rect 3965 5956 3989 5958
rect 4045 5956 4069 5958
rect 4125 5956 4131 5958
rect 3823 5947 4131 5956
rect 5800 6012 6108 6021
rect 5800 6010 5806 6012
rect 5862 6010 5886 6012
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6108 6012
rect 5862 5958 5864 6010
rect 6044 5958 6046 6010
rect 5800 5956 5806 5958
rect 5862 5956 5886 5958
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6108 5958
rect 5800 5947 6108 5956
rect 7777 6012 8085 6021
rect 7777 6010 7783 6012
rect 7839 6010 7863 6012
rect 7919 6010 7943 6012
rect 7999 6010 8023 6012
rect 8079 6010 8085 6012
rect 7839 5958 7841 6010
rect 8021 5958 8023 6010
rect 7777 5956 7783 5958
rect 7839 5956 7863 5958
rect 7919 5956 7943 5958
rect 7999 5956 8023 5958
rect 8079 5956 8085 5958
rect 7777 5947 8085 5956
rect 2834 5468 3142 5477
rect 2834 5466 2840 5468
rect 2896 5466 2920 5468
rect 2976 5466 3000 5468
rect 3056 5466 3080 5468
rect 3136 5466 3142 5468
rect 2896 5414 2898 5466
rect 3078 5414 3080 5466
rect 2834 5412 2840 5414
rect 2896 5412 2920 5414
rect 2976 5412 3000 5414
rect 3056 5412 3080 5414
rect 3136 5412 3142 5414
rect 2834 5403 3142 5412
rect 4811 5468 5119 5477
rect 4811 5466 4817 5468
rect 4873 5466 4897 5468
rect 4953 5466 4977 5468
rect 5033 5466 5057 5468
rect 5113 5466 5119 5468
rect 4873 5414 4875 5466
rect 5055 5414 5057 5466
rect 4811 5412 4817 5414
rect 4873 5412 4897 5414
rect 4953 5412 4977 5414
rect 5033 5412 5057 5414
rect 5113 5412 5119 5414
rect 4811 5403 5119 5412
rect 6788 5468 7096 5477
rect 6788 5466 6794 5468
rect 6850 5466 6874 5468
rect 6930 5466 6954 5468
rect 7010 5466 7034 5468
rect 7090 5466 7096 5468
rect 6850 5414 6852 5466
rect 7032 5414 7034 5466
rect 6788 5412 6794 5414
rect 6850 5412 6874 5414
rect 6930 5412 6954 5414
rect 7010 5412 7034 5414
rect 7090 5412 7096 5414
rect 6788 5403 7096 5412
rect 8312 5098 8340 6734
rect 8404 5302 8432 6734
rect 8765 6556 9073 6565
rect 8765 6554 8771 6556
rect 8827 6554 8851 6556
rect 8907 6554 8931 6556
rect 8987 6554 9011 6556
rect 9067 6554 9073 6556
rect 8827 6502 8829 6554
rect 9009 6502 9011 6554
rect 8765 6500 8771 6502
rect 8827 6500 8851 6502
rect 8907 6500 8931 6502
rect 8987 6500 9011 6502
rect 9067 6500 9073 6502
rect 8765 6491 9073 6500
rect 8765 5468 9073 5477
rect 8765 5466 8771 5468
rect 8827 5466 8851 5468
rect 8907 5466 8931 5468
rect 8987 5466 9011 5468
rect 9067 5466 9073 5468
rect 8827 5414 8829 5466
rect 9009 5414 9011 5466
rect 8765 5412 8771 5414
rect 8827 5412 8851 5414
rect 8907 5412 8931 5414
rect 8987 5412 9011 5414
rect 9067 5412 9073 5414
rect 8765 5403 9073 5412
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8208 5024 8260 5030
rect 8206 4992 8208 5001
rect 8260 4992 8262 5001
rect 1846 4924 2154 4933
rect 1846 4922 1852 4924
rect 1908 4922 1932 4924
rect 1988 4922 2012 4924
rect 2068 4922 2092 4924
rect 2148 4922 2154 4924
rect 1908 4870 1910 4922
rect 2090 4870 2092 4922
rect 1846 4868 1852 4870
rect 1908 4868 1932 4870
rect 1988 4868 2012 4870
rect 2068 4868 2092 4870
rect 2148 4868 2154 4870
rect 1846 4859 2154 4868
rect 3823 4924 4131 4933
rect 3823 4922 3829 4924
rect 3885 4922 3909 4924
rect 3965 4922 3989 4924
rect 4045 4922 4069 4924
rect 4125 4922 4131 4924
rect 3885 4870 3887 4922
rect 4067 4870 4069 4922
rect 3823 4868 3829 4870
rect 3885 4868 3909 4870
rect 3965 4868 3989 4870
rect 4045 4868 4069 4870
rect 4125 4868 4131 4870
rect 3823 4859 4131 4868
rect 5800 4924 6108 4933
rect 5800 4922 5806 4924
rect 5862 4922 5886 4924
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6108 4924
rect 5862 4870 5864 4922
rect 6044 4870 6046 4922
rect 5800 4868 5806 4870
rect 5862 4868 5886 4870
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6108 4870
rect 5800 4859 6108 4868
rect 7777 4924 8085 4933
rect 8206 4927 8262 4936
rect 7777 4922 7783 4924
rect 7839 4922 7863 4924
rect 7919 4922 7943 4924
rect 7999 4922 8023 4924
rect 8079 4922 8085 4924
rect 7839 4870 7841 4922
rect 8021 4870 8023 4922
rect 7777 4868 7783 4870
rect 7839 4868 7863 4870
rect 7919 4868 7943 4870
rect 7999 4868 8023 4870
rect 8079 4868 8085 4870
rect 7777 4859 8085 4868
rect 2834 4380 3142 4389
rect 2834 4378 2840 4380
rect 2896 4378 2920 4380
rect 2976 4378 3000 4380
rect 3056 4378 3080 4380
rect 3136 4378 3142 4380
rect 2896 4326 2898 4378
rect 3078 4326 3080 4378
rect 2834 4324 2840 4326
rect 2896 4324 2920 4326
rect 2976 4324 3000 4326
rect 3056 4324 3080 4326
rect 3136 4324 3142 4326
rect 2834 4315 3142 4324
rect 4811 4380 5119 4389
rect 4811 4378 4817 4380
rect 4873 4378 4897 4380
rect 4953 4378 4977 4380
rect 5033 4378 5057 4380
rect 5113 4378 5119 4380
rect 4873 4326 4875 4378
rect 5055 4326 5057 4378
rect 4811 4324 4817 4326
rect 4873 4324 4897 4326
rect 4953 4324 4977 4326
rect 5033 4324 5057 4326
rect 5113 4324 5119 4326
rect 4811 4315 5119 4324
rect 6788 4380 7096 4389
rect 6788 4378 6794 4380
rect 6850 4378 6874 4380
rect 6930 4378 6954 4380
rect 7010 4378 7034 4380
rect 7090 4378 7096 4380
rect 6850 4326 6852 4378
rect 7032 4326 7034 4378
rect 6788 4324 6794 4326
rect 6850 4324 6874 4326
rect 6930 4324 6954 4326
rect 7010 4324 7034 4326
rect 7090 4324 7096 4326
rect 6788 4315 7096 4324
rect 1846 3836 2154 3845
rect 1846 3834 1852 3836
rect 1908 3834 1932 3836
rect 1988 3834 2012 3836
rect 2068 3834 2092 3836
rect 2148 3834 2154 3836
rect 1908 3782 1910 3834
rect 2090 3782 2092 3834
rect 1846 3780 1852 3782
rect 1908 3780 1932 3782
rect 1988 3780 2012 3782
rect 2068 3780 2092 3782
rect 2148 3780 2154 3782
rect 1846 3771 2154 3780
rect 3823 3836 4131 3845
rect 3823 3834 3829 3836
rect 3885 3834 3909 3836
rect 3965 3834 3989 3836
rect 4045 3834 4069 3836
rect 4125 3834 4131 3836
rect 3885 3782 3887 3834
rect 4067 3782 4069 3834
rect 3823 3780 3829 3782
rect 3885 3780 3909 3782
rect 3965 3780 3989 3782
rect 4045 3780 4069 3782
rect 4125 3780 4131 3782
rect 3823 3771 4131 3780
rect 5800 3836 6108 3845
rect 5800 3834 5806 3836
rect 5862 3834 5886 3836
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6108 3836
rect 5862 3782 5864 3834
rect 6044 3782 6046 3834
rect 5800 3780 5806 3782
rect 5862 3780 5886 3782
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6108 3782
rect 5800 3771 6108 3780
rect 7777 3836 8085 3845
rect 7777 3834 7783 3836
rect 7839 3834 7863 3836
rect 7919 3834 7943 3836
rect 7999 3834 8023 3836
rect 8079 3834 8085 3836
rect 7839 3782 7841 3834
rect 8021 3782 8023 3834
rect 7777 3780 7783 3782
rect 7839 3780 7863 3782
rect 7919 3780 7943 3782
rect 7999 3780 8023 3782
rect 8079 3780 8085 3782
rect 7777 3771 8085 3780
rect 2834 3292 3142 3301
rect 2834 3290 2840 3292
rect 2896 3290 2920 3292
rect 2976 3290 3000 3292
rect 3056 3290 3080 3292
rect 3136 3290 3142 3292
rect 2896 3238 2898 3290
rect 3078 3238 3080 3290
rect 2834 3236 2840 3238
rect 2896 3236 2920 3238
rect 2976 3236 3000 3238
rect 3056 3236 3080 3238
rect 3136 3236 3142 3238
rect 2834 3227 3142 3236
rect 4811 3292 5119 3301
rect 4811 3290 4817 3292
rect 4873 3290 4897 3292
rect 4953 3290 4977 3292
rect 5033 3290 5057 3292
rect 5113 3290 5119 3292
rect 4873 3238 4875 3290
rect 5055 3238 5057 3290
rect 4811 3236 4817 3238
rect 4873 3236 4897 3238
rect 4953 3236 4977 3238
rect 5033 3236 5057 3238
rect 5113 3236 5119 3238
rect 4811 3227 5119 3236
rect 6788 3292 7096 3301
rect 6788 3290 6794 3292
rect 6850 3290 6874 3292
rect 6930 3290 6954 3292
rect 7010 3290 7034 3292
rect 7090 3290 7096 3292
rect 6850 3238 6852 3290
rect 7032 3238 7034 3290
rect 6788 3236 6794 3238
rect 6850 3236 6874 3238
rect 6930 3236 6954 3238
rect 7010 3236 7034 3238
rect 7090 3236 7096 3238
rect 6788 3227 7096 3236
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7668 3097 7696 3130
rect 7654 3088 7710 3097
rect 8312 3058 8340 5034
rect 7654 3023 7710 3032
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8404 2938 8432 5238
rect 8765 4380 9073 4389
rect 8765 4378 8771 4380
rect 8827 4378 8851 4380
rect 8907 4378 8931 4380
rect 8987 4378 9011 4380
rect 9067 4378 9073 4380
rect 8827 4326 8829 4378
rect 9009 4326 9011 4378
rect 8765 4324 8771 4326
rect 8827 4324 8851 4326
rect 8907 4324 8931 4326
rect 8987 4324 9011 4326
rect 9067 4324 9073 4326
rect 8765 4315 9073 4324
rect 8765 3292 9073 3301
rect 8765 3290 8771 3292
rect 8827 3290 8851 3292
rect 8907 3290 8931 3292
rect 8987 3290 9011 3292
rect 9067 3290 9073 3292
rect 8827 3238 8829 3290
rect 9009 3238 9011 3290
rect 8765 3236 8771 3238
rect 8827 3236 8851 3238
rect 8907 3236 8931 3238
rect 8987 3236 9011 3238
rect 9067 3236 9073 3238
rect 8765 3227 9073 3236
rect 8312 2922 8432 2938
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8300 2916 8432 2922
rect 8352 2910 8432 2916
rect 8300 2858 8352 2864
rect 1846 2748 2154 2757
rect 1846 2746 1852 2748
rect 1908 2746 1932 2748
rect 1988 2746 2012 2748
rect 2068 2746 2092 2748
rect 2148 2746 2154 2748
rect 1908 2694 1910 2746
rect 2090 2694 2092 2746
rect 1846 2692 1852 2694
rect 1908 2692 1932 2694
rect 1988 2692 2012 2694
rect 2068 2692 2092 2694
rect 2148 2692 2154 2694
rect 1846 2683 2154 2692
rect 3823 2748 4131 2757
rect 3823 2746 3829 2748
rect 3885 2746 3909 2748
rect 3965 2746 3989 2748
rect 4045 2746 4069 2748
rect 4125 2746 4131 2748
rect 3885 2694 3887 2746
rect 4067 2694 4069 2746
rect 3823 2692 3829 2694
rect 3885 2692 3909 2694
rect 3965 2692 3989 2694
rect 4045 2692 4069 2694
rect 4125 2692 4131 2694
rect 3823 2683 4131 2692
rect 5800 2748 6108 2757
rect 5800 2746 5806 2748
rect 5862 2746 5886 2748
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6108 2748
rect 5862 2694 5864 2746
rect 6044 2694 6046 2746
rect 5800 2692 5806 2694
rect 5862 2692 5886 2694
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6108 2694
rect 5800 2683 6108 2692
rect 7777 2748 8085 2757
rect 7777 2746 7783 2748
rect 7839 2746 7863 2748
rect 7919 2746 7943 2748
rect 7999 2746 8023 2748
rect 8079 2746 8085 2748
rect 7839 2694 7841 2746
rect 8021 2694 8023 2746
rect 7777 2692 7783 2694
rect 7839 2692 7863 2694
rect 7919 2692 7943 2694
rect 7999 2692 8023 2694
rect 8079 2692 8085 2694
rect 7777 2683 8085 2692
rect 2834 2204 3142 2213
rect 2834 2202 2840 2204
rect 2896 2202 2920 2204
rect 2976 2202 3000 2204
rect 3056 2202 3080 2204
rect 3136 2202 3142 2204
rect 2896 2150 2898 2202
rect 3078 2150 3080 2202
rect 2834 2148 2840 2150
rect 2896 2148 2920 2150
rect 2976 2148 3000 2150
rect 3056 2148 3080 2150
rect 3136 2148 3142 2150
rect 2834 2139 3142 2148
rect 4811 2204 5119 2213
rect 4811 2202 4817 2204
rect 4873 2202 4897 2204
rect 4953 2202 4977 2204
rect 5033 2202 5057 2204
rect 5113 2202 5119 2204
rect 4873 2150 4875 2202
rect 5055 2150 5057 2202
rect 4811 2148 4817 2150
rect 4873 2148 4897 2150
rect 4953 2148 4977 2150
rect 5033 2148 5057 2150
rect 5113 2148 5119 2150
rect 4811 2139 5119 2148
rect 6788 2204 7096 2213
rect 6788 2202 6794 2204
rect 6850 2202 6874 2204
rect 6930 2202 6954 2204
rect 7010 2202 7034 2204
rect 7090 2202 7096 2204
rect 6850 2150 6852 2202
rect 7032 2150 7034 2202
rect 6788 2148 6794 2150
rect 6850 2148 6874 2150
rect 6930 2148 6954 2150
rect 7010 2148 7034 2150
rect 7090 2148 7096 2150
rect 6788 2139 7096 2148
rect 8128 1970 8156 2858
rect 8392 2848 8444 2854
rect 8312 2796 8392 2802
rect 8312 2790 8444 2796
rect 8312 2774 8432 2790
rect 8312 1970 8340 2774
rect 8765 2204 9073 2213
rect 8765 2202 8771 2204
rect 8827 2202 8851 2204
rect 8907 2202 8931 2204
rect 8987 2202 9011 2204
rect 9067 2202 9073 2204
rect 8827 2150 8829 2202
rect 9009 2150 9011 2202
rect 8765 2148 8771 2150
rect 8827 2148 8851 2150
rect 8907 2148 8931 2150
rect 8987 2148 9011 2150
rect 9067 2148 9073 2150
rect 8765 2139 9073 2148
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 1846 1660 2154 1669
rect 1846 1658 1852 1660
rect 1908 1658 1932 1660
rect 1988 1658 2012 1660
rect 2068 1658 2092 1660
rect 2148 1658 2154 1660
rect 1908 1606 1910 1658
rect 2090 1606 2092 1658
rect 1846 1604 1852 1606
rect 1908 1604 1932 1606
rect 1988 1604 2012 1606
rect 2068 1604 2092 1606
rect 2148 1604 2154 1606
rect 1846 1595 2154 1604
rect 3823 1660 4131 1669
rect 3823 1658 3829 1660
rect 3885 1658 3909 1660
rect 3965 1658 3989 1660
rect 4045 1658 4069 1660
rect 4125 1658 4131 1660
rect 3885 1606 3887 1658
rect 4067 1606 4069 1658
rect 3823 1604 3829 1606
rect 3885 1604 3909 1606
rect 3965 1604 3989 1606
rect 4045 1604 4069 1606
rect 4125 1604 4131 1606
rect 3823 1595 4131 1604
rect 5800 1660 6108 1669
rect 5800 1658 5806 1660
rect 5862 1658 5886 1660
rect 5942 1658 5966 1660
rect 6022 1658 6046 1660
rect 6102 1658 6108 1660
rect 5862 1606 5864 1658
rect 6044 1606 6046 1658
rect 5800 1604 5806 1606
rect 5862 1604 5886 1606
rect 5942 1604 5966 1606
rect 6022 1604 6046 1606
rect 6102 1604 6108 1606
rect 5800 1595 6108 1604
rect 7777 1660 8085 1669
rect 7777 1658 7783 1660
rect 7839 1658 7863 1660
rect 7919 1658 7943 1660
rect 7999 1658 8023 1660
rect 8079 1658 8085 1660
rect 7839 1606 7841 1658
rect 8021 1606 8023 1658
rect 7777 1604 7783 1606
rect 7839 1604 7863 1606
rect 7919 1604 7943 1606
rect 7999 1604 8023 1606
rect 8079 1604 8085 1606
rect 7777 1595 8085 1604
rect 8128 1562 8156 1906
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8312 1494 8340 1906
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 8300 1488 8352 1494
rect 8300 1430 8352 1436
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 2504 1284 2556 1290
rect 2504 1226 2556 1232
rect 2516 400 2544 1226
rect 2834 1116 3142 1125
rect 2834 1114 2840 1116
rect 2896 1114 2920 1116
rect 2976 1114 3000 1116
rect 3056 1114 3080 1116
rect 3136 1114 3142 1116
rect 2896 1062 2898 1114
rect 3078 1062 3080 1114
rect 2834 1060 2840 1062
rect 2896 1060 2920 1062
rect 2976 1060 3000 1062
rect 3056 1060 3080 1062
rect 3136 1060 3142 1062
rect 2834 1051 3142 1060
rect 4811 1116 5119 1125
rect 4811 1114 4817 1116
rect 4873 1114 4897 1116
rect 4953 1114 4977 1116
rect 5033 1114 5057 1116
rect 5113 1114 5119 1116
rect 4873 1062 4875 1114
rect 5055 1062 5057 1114
rect 4811 1060 4817 1062
rect 4873 1060 4897 1062
rect 4953 1060 4977 1062
rect 5033 1060 5057 1062
rect 5113 1060 5119 1062
rect 4811 1051 5119 1060
rect 6788 1116 7096 1125
rect 6788 1114 6794 1116
rect 6850 1114 6874 1116
rect 6930 1114 6954 1116
rect 7010 1114 7034 1116
rect 7090 1114 7096 1116
rect 6850 1062 6852 1114
rect 7032 1062 7034 1114
rect 6788 1060 6794 1062
rect 6850 1060 6874 1062
rect 6930 1060 6954 1062
rect 7010 1060 7034 1062
rect 7090 1060 7096 1062
rect 6788 1051 7096 1060
rect 7484 400 7512 1294
rect 9324 1193 9352 1838
rect 9310 1184 9366 1193
rect 8765 1116 9073 1125
rect 9310 1119 9366 1128
rect 8765 1114 8771 1116
rect 8827 1114 8851 1116
rect 8907 1114 8931 1116
rect 8987 1114 9011 1116
rect 9067 1114 9073 1116
rect 8827 1062 8829 1114
rect 9009 1062 9011 1114
rect 8765 1060 8771 1062
rect 8827 1060 8851 1062
rect 8907 1060 8931 1062
rect 8987 1060 9011 1062
rect 9067 1060 9073 1062
rect 8765 1051 9073 1060
rect 2502 0 2558 400
rect 7470 0 7526 400
<< via2 >>
rect 1852 14714 1908 14716
rect 1932 14714 1988 14716
rect 2012 14714 2068 14716
rect 2092 14714 2148 14716
rect 1852 14662 1898 14714
rect 1898 14662 1908 14714
rect 1932 14662 1962 14714
rect 1962 14662 1974 14714
rect 1974 14662 1988 14714
rect 2012 14662 2026 14714
rect 2026 14662 2038 14714
rect 2038 14662 2068 14714
rect 2092 14662 2102 14714
rect 2102 14662 2148 14714
rect 1852 14660 1908 14662
rect 1932 14660 1988 14662
rect 2012 14660 2068 14662
rect 2092 14660 2148 14662
rect 3829 14714 3885 14716
rect 3909 14714 3965 14716
rect 3989 14714 4045 14716
rect 4069 14714 4125 14716
rect 3829 14662 3875 14714
rect 3875 14662 3885 14714
rect 3909 14662 3939 14714
rect 3939 14662 3951 14714
rect 3951 14662 3965 14714
rect 3989 14662 4003 14714
rect 4003 14662 4015 14714
rect 4015 14662 4045 14714
rect 4069 14662 4079 14714
rect 4079 14662 4125 14714
rect 3829 14660 3885 14662
rect 3909 14660 3965 14662
rect 3989 14660 4045 14662
rect 4069 14660 4125 14662
rect 5806 14714 5862 14716
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 5806 14662 5852 14714
rect 5852 14662 5862 14714
rect 5886 14662 5916 14714
rect 5916 14662 5928 14714
rect 5928 14662 5942 14714
rect 5966 14662 5980 14714
rect 5980 14662 5992 14714
rect 5992 14662 6022 14714
rect 6046 14662 6056 14714
rect 6056 14662 6102 14714
rect 5806 14660 5862 14662
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 7783 14714 7839 14716
rect 7863 14714 7919 14716
rect 7943 14714 7999 14716
rect 8023 14714 8079 14716
rect 7783 14662 7829 14714
rect 7829 14662 7839 14714
rect 7863 14662 7893 14714
rect 7893 14662 7905 14714
rect 7905 14662 7919 14714
rect 7943 14662 7957 14714
rect 7957 14662 7969 14714
rect 7969 14662 7999 14714
rect 8023 14662 8033 14714
rect 8033 14662 8079 14714
rect 7783 14660 7839 14662
rect 7863 14660 7919 14662
rect 7943 14660 7999 14662
rect 8023 14660 8079 14662
rect 8114 14456 8170 14512
rect 2840 14170 2896 14172
rect 2920 14170 2976 14172
rect 3000 14170 3056 14172
rect 3080 14170 3136 14172
rect 2840 14118 2886 14170
rect 2886 14118 2896 14170
rect 2920 14118 2950 14170
rect 2950 14118 2962 14170
rect 2962 14118 2976 14170
rect 3000 14118 3014 14170
rect 3014 14118 3026 14170
rect 3026 14118 3056 14170
rect 3080 14118 3090 14170
rect 3090 14118 3136 14170
rect 2840 14116 2896 14118
rect 2920 14116 2976 14118
rect 3000 14116 3056 14118
rect 3080 14116 3136 14118
rect 4817 14170 4873 14172
rect 4897 14170 4953 14172
rect 4977 14170 5033 14172
rect 5057 14170 5113 14172
rect 4817 14118 4863 14170
rect 4863 14118 4873 14170
rect 4897 14118 4927 14170
rect 4927 14118 4939 14170
rect 4939 14118 4953 14170
rect 4977 14118 4991 14170
rect 4991 14118 5003 14170
rect 5003 14118 5033 14170
rect 5057 14118 5067 14170
rect 5067 14118 5113 14170
rect 4817 14116 4873 14118
rect 4897 14116 4953 14118
rect 4977 14116 5033 14118
rect 5057 14116 5113 14118
rect 6794 14170 6850 14172
rect 6874 14170 6930 14172
rect 6954 14170 7010 14172
rect 7034 14170 7090 14172
rect 6794 14118 6840 14170
rect 6840 14118 6850 14170
rect 6874 14118 6904 14170
rect 6904 14118 6916 14170
rect 6916 14118 6930 14170
rect 6954 14118 6968 14170
rect 6968 14118 6980 14170
rect 6980 14118 7010 14170
rect 7034 14118 7044 14170
rect 7044 14118 7090 14170
rect 6794 14116 6850 14118
rect 6874 14116 6930 14118
rect 6954 14116 7010 14118
rect 7034 14116 7090 14118
rect 1852 13626 1908 13628
rect 1932 13626 1988 13628
rect 2012 13626 2068 13628
rect 2092 13626 2148 13628
rect 1852 13574 1898 13626
rect 1898 13574 1908 13626
rect 1932 13574 1962 13626
rect 1962 13574 1974 13626
rect 1974 13574 1988 13626
rect 2012 13574 2026 13626
rect 2026 13574 2038 13626
rect 2038 13574 2068 13626
rect 2092 13574 2102 13626
rect 2102 13574 2148 13626
rect 1852 13572 1908 13574
rect 1932 13572 1988 13574
rect 2012 13572 2068 13574
rect 2092 13572 2148 13574
rect 3829 13626 3885 13628
rect 3909 13626 3965 13628
rect 3989 13626 4045 13628
rect 4069 13626 4125 13628
rect 3829 13574 3875 13626
rect 3875 13574 3885 13626
rect 3909 13574 3939 13626
rect 3939 13574 3951 13626
rect 3951 13574 3965 13626
rect 3989 13574 4003 13626
rect 4003 13574 4015 13626
rect 4015 13574 4045 13626
rect 4069 13574 4079 13626
rect 4079 13574 4125 13626
rect 3829 13572 3885 13574
rect 3909 13572 3965 13574
rect 3989 13572 4045 13574
rect 4069 13572 4125 13574
rect 5806 13626 5862 13628
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 5806 13574 5852 13626
rect 5852 13574 5862 13626
rect 5886 13574 5916 13626
rect 5916 13574 5928 13626
rect 5928 13574 5942 13626
rect 5966 13574 5980 13626
rect 5980 13574 5992 13626
rect 5992 13574 6022 13626
rect 6046 13574 6056 13626
rect 6056 13574 6102 13626
rect 5806 13572 5862 13574
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 7783 13626 7839 13628
rect 7863 13626 7919 13628
rect 7943 13626 7999 13628
rect 8023 13626 8079 13628
rect 7783 13574 7829 13626
rect 7829 13574 7839 13626
rect 7863 13574 7893 13626
rect 7893 13574 7905 13626
rect 7905 13574 7919 13626
rect 7943 13574 7957 13626
rect 7957 13574 7969 13626
rect 7969 13574 7999 13626
rect 8023 13574 8033 13626
rect 8033 13574 8079 13626
rect 7783 13572 7839 13574
rect 7863 13572 7919 13574
rect 7943 13572 7999 13574
rect 8023 13572 8079 13574
rect 2840 13082 2896 13084
rect 2920 13082 2976 13084
rect 3000 13082 3056 13084
rect 3080 13082 3136 13084
rect 2840 13030 2886 13082
rect 2886 13030 2896 13082
rect 2920 13030 2950 13082
rect 2950 13030 2962 13082
rect 2962 13030 2976 13082
rect 3000 13030 3014 13082
rect 3014 13030 3026 13082
rect 3026 13030 3056 13082
rect 3080 13030 3090 13082
rect 3090 13030 3136 13082
rect 2840 13028 2896 13030
rect 2920 13028 2976 13030
rect 3000 13028 3056 13030
rect 3080 13028 3136 13030
rect 4817 13082 4873 13084
rect 4897 13082 4953 13084
rect 4977 13082 5033 13084
rect 5057 13082 5113 13084
rect 4817 13030 4863 13082
rect 4863 13030 4873 13082
rect 4897 13030 4927 13082
rect 4927 13030 4939 13082
rect 4939 13030 4953 13082
rect 4977 13030 4991 13082
rect 4991 13030 5003 13082
rect 5003 13030 5033 13082
rect 5057 13030 5067 13082
rect 5067 13030 5113 13082
rect 4817 13028 4873 13030
rect 4897 13028 4953 13030
rect 4977 13028 5033 13030
rect 5057 13028 5113 13030
rect 6794 13082 6850 13084
rect 6874 13082 6930 13084
rect 6954 13082 7010 13084
rect 7034 13082 7090 13084
rect 6794 13030 6840 13082
rect 6840 13030 6850 13082
rect 6874 13030 6904 13082
rect 6904 13030 6916 13082
rect 6916 13030 6930 13082
rect 6954 13030 6968 13082
rect 6968 13030 6980 13082
rect 6980 13030 7010 13082
rect 7034 13030 7044 13082
rect 7044 13030 7090 13082
rect 6794 13028 6850 13030
rect 6874 13028 6930 13030
rect 6954 13028 7010 13030
rect 7034 13028 7090 13030
rect 1852 12538 1908 12540
rect 1932 12538 1988 12540
rect 2012 12538 2068 12540
rect 2092 12538 2148 12540
rect 1852 12486 1898 12538
rect 1898 12486 1908 12538
rect 1932 12486 1962 12538
rect 1962 12486 1974 12538
rect 1974 12486 1988 12538
rect 2012 12486 2026 12538
rect 2026 12486 2038 12538
rect 2038 12486 2068 12538
rect 2092 12486 2102 12538
rect 2102 12486 2148 12538
rect 1852 12484 1908 12486
rect 1932 12484 1988 12486
rect 2012 12484 2068 12486
rect 2092 12484 2148 12486
rect 3829 12538 3885 12540
rect 3909 12538 3965 12540
rect 3989 12538 4045 12540
rect 4069 12538 4125 12540
rect 3829 12486 3875 12538
rect 3875 12486 3885 12538
rect 3909 12486 3939 12538
rect 3939 12486 3951 12538
rect 3951 12486 3965 12538
rect 3989 12486 4003 12538
rect 4003 12486 4015 12538
rect 4015 12486 4045 12538
rect 4069 12486 4079 12538
rect 4079 12486 4125 12538
rect 3829 12484 3885 12486
rect 3909 12484 3965 12486
rect 3989 12484 4045 12486
rect 4069 12484 4125 12486
rect 5806 12538 5862 12540
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 5806 12486 5852 12538
rect 5852 12486 5862 12538
rect 5886 12486 5916 12538
rect 5916 12486 5928 12538
rect 5928 12486 5942 12538
rect 5966 12486 5980 12538
rect 5980 12486 5992 12538
rect 5992 12486 6022 12538
rect 6046 12486 6056 12538
rect 6056 12486 6102 12538
rect 5806 12484 5862 12486
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 7783 12538 7839 12540
rect 7863 12538 7919 12540
rect 7943 12538 7999 12540
rect 8023 12538 8079 12540
rect 7783 12486 7829 12538
rect 7829 12486 7839 12538
rect 7863 12486 7893 12538
rect 7893 12486 7905 12538
rect 7905 12486 7919 12538
rect 7943 12486 7957 12538
rect 7957 12486 7969 12538
rect 7969 12486 7999 12538
rect 8023 12486 8033 12538
rect 8033 12486 8079 12538
rect 7783 12484 7839 12486
rect 7863 12484 7919 12486
rect 7943 12484 7999 12486
rect 8023 12484 8079 12486
rect 2840 11994 2896 11996
rect 2920 11994 2976 11996
rect 3000 11994 3056 11996
rect 3080 11994 3136 11996
rect 2840 11942 2886 11994
rect 2886 11942 2896 11994
rect 2920 11942 2950 11994
rect 2950 11942 2962 11994
rect 2962 11942 2976 11994
rect 3000 11942 3014 11994
rect 3014 11942 3026 11994
rect 3026 11942 3056 11994
rect 3080 11942 3090 11994
rect 3090 11942 3136 11994
rect 2840 11940 2896 11942
rect 2920 11940 2976 11942
rect 3000 11940 3056 11942
rect 3080 11940 3136 11942
rect 4817 11994 4873 11996
rect 4897 11994 4953 11996
rect 4977 11994 5033 11996
rect 5057 11994 5113 11996
rect 4817 11942 4863 11994
rect 4863 11942 4873 11994
rect 4897 11942 4927 11994
rect 4927 11942 4939 11994
rect 4939 11942 4953 11994
rect 4977 11942 4991 11994
rect 4991 11942 5003 11994
rect 5003 11942 5033 11994
rect 5057 11942 5067 11994
rect 5067 11942 5113 11994
rect 4817 11940 4873 11942
rect 4897 11940 4953 11942
rect 4977 11940 5033 11942
rect 5057 11940 5113 11942
rect 6794 11994 6850 11996
rect 6874 11994 6930 11996
rect 6954 11994 7010 11996
rect 7034 11994 7090 11996
rect 6794 11942 6840 11994
rect 6840 11942 6850 11994
rect 6874 11942 6904 11994
rect 6904 11942 6916 11994
rect 6916 11942 6930 11994
rect 6954 11942 6968 11994
rect 6968 11942 6980 11994
rect 6980 11942 7010 11994
rect 7034 11942 7044 11994
rect 7044 11942 7090 11994
rect 6794 11940 6850 11942
rect 6874 11940 6930 11942
rect 6954 11940 7010 11942
rect 7034 11940 7090 11942
rect 8771 14170 8827 14172
rect 8851 14170 8907 14172
rect 8931 14170 8987 14172
rect 9011 14170 9067 14172
rect 8771 14118 8817 14170
rect 8817 14118 8827 14170
rect 8851 14118 8881 14170
rect 8881 14118 8893 14170
rect 8893 14118 8907 14170
rect 8931 14118 8945 14170
rect 8945 14118 8957 14170
rect 8957 14118 8987 14170
rect 9011 14118 9021 14170
rect 9021 14118 9067 14170
rect 8771 14116 8827 14118
rect 8851 14116 8907 14118
rect 8931 14116 8987 14118
rect 9011 14116 9067 14118
rect 8771 13082 8827 13084
rect 8851 13082 8907 13084
rect 8931 13082 8987 13084
rect 9011 13082 9067 13084
rect 8771 13030 8817 13082
rect 8817 13030 8827 13082
rect 8851 13030 8881 13082
rect 8881 13030 8893 13082
rect 8893 13030 8907 13082
rect 8931 13030 8945 13082
rect 8945 13030 8957 13082
rect 8957 13030 8987 13082
rect 9011 13030 9021 13082
rect 9021 13030 9067 13082
rect 8771 13028 8827 13030
rect 8851 13028 8907 13030
rect 8931 13028 8987 13030
rect 9011 13028 9067 13030
rect 8206 12552 8262 12608
rect 1852 11450 1908 11452
rect 1932 11450 1988 11452
rect 2012 11450 2068 11452
rect 2092 11450 2148 11452
rect 1852 11398 1898 11450
rect 1898 11398 1908 11450
rect 1932 11398 1962 11450
rect 1962 11398 1974 11450
rect 1974 11398 1988 11450
rect 2012 11398 2026 11450
rect 2026 11398 2038 11450
rect 2038 11398 2068 11450
rect 2092 11398 2102 11450
rect 2102 11398 2148 11450
rect 1852 11396 1908 11398
rect 1932 11396 1988 11398
rect 2012 11396 2068 11398
rect 2092 11396 2148 11398
rect 3829 11450 3885 11452
rect 3909 11450 3965 11452
rect 3989 11450 4045 11452
rect 4069 11450 4125 11452
rect 3829 11398 3875 11450
rect 3875 11398 3885 11450
rect 3909 11398 3939 11450
rect 3939 11398 3951 11450
rect 3951 11398 3965 11450
rect 3989 11398 4003 11450
rect 4003 11398 4015 11450
rect 4015 11398 4045 11450
rect 4069 11398 4079 11450
rect 4079 11398 4125 11450
rect 3829 11396 3885 11398
rect 3909 11396 3965 11398
rect 3989 11396 4045 11398
rect 4069 11396 4125 11398
rect 5806 11450 5862 11452
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 5806 11398 5852 11450
rect 5852 11398 5862 11450
rect 5886 11398 5916 11450
rect 5916 11398 5928 11450
rect 5928 11398 5942 11450
rect 5966 11398 5980 11450
rect 5980 11398 5992 11450
rect 5992 11398 6022 11450
rect 6046 11398 6056 11450
rect 6056 11398 6102 11450
rect 5806 11396 5862 11398
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 7783 11450 7839 11452
rect 7863 11450 7919 11452
rect 7943 11450 7999 11452
rect 8023 11450 8079 11452
rect 7783 11398 7829 11450
rect 7829 11398 7839 11450
rect 7863 11398 7893 11450
rect 7893 11398 7905 11450
rect 7905 11398 7919 11450
rect 7943 11398 7957 11450
rect 7957 11398 7969 11450
rect 7969 11398 7999 11450
rect 8023 11398 8033 11450
rect 8033 11398 8079 11450
rect 7783 11396 7839 11398
rect 7863 11396 7919 11398
rect 7943 11396 7999 11398
rect 8023 11396 8079 11398
rect 8771 11994 8827 11996
rect 8851 11994 8907 11996
rect 8931 11994 8987 11996
rect 9011 11994 9067 11996
rect 8771 11942 8817 11994
rect 8817 11942 8827 11994
rect 8851 11942 8881 11994
rect 8881 11942 8893 11994
rect 8893 11942 8907 11994
rect 8931 11942 8945 11994
rect 8945 11942 8957 11994
rect 8957 11942 8987 11994
rect 9011 11942 9021 11994
rect 9021 11942 9067 11994
rect 8771 11940 8827 11942
rect 8851 11940 8907 11942
rect 8931 11940 8987 11942
rect 9011 11940 9067 11942
rect 2840 10906 2896 10908
rect 2920 10906 2976 10908
rect 3000 10906 3056 10908
rect 3080 10906 3136 10908
rect 2840 10854 2886 10906
rect 2886 10854 2896 10906
rect 2920 10854 2950 10906
rect 2950 10854 2962 10906
rect 2962 10854 2976 10906
rect 3000 10854 3014 10906
rect 3014 10854 3026 10906
rect 3026 10854 3056 10906
rect 3080 10854 3090 10906
rect 3090 10854 3136 10906
rect 2840 10852 2896 10854
rect 2920 10852 2976 10854
rect 3000 10852 3056 10854
rect 3080 10852 3136 10854
rect 4817 10906 4873 10908
rect 4897 10906 4953 10908
rect 4977 10906 5033 10908
rect 5057 10906 5113 10908
rect 4817 10854 4863 10906
rect 4863 10854 4873 10906
rect 4897 10854 4927 10906
rect 4927 10854 4939 10906
rect 4939 10854 4953 10906
rect 4977 10854 4991 10906
rect 4991 10854 5003 10906
rect 5003 10854 5033 10906
rect 5057 10854 5067 10906
rect 5067 10854 5113 10906
rect 4817 10852 4873 10854
rect 4897 10852 4953 10854
rect 4977 10852 5033 10854
rect 5057 10852 5113 10854
rect 6794 10906 6850 10908
rect 6874 10906 6930 10908
rect 6954 10906 7010 10908
rect 7034 10906 7090 10908
rect 6794 10854 6840 10906
rect 6840 10854 6850 10906
rect 6874 10854 6904 10906
rect 6904 10854 6916 10906
rect 6916 10854 6930 10906
rect 6954 10854 6968 10906
rect 6968 10854 6980 10906
rect 6980 10854 7010 10906
rect 7034 10854 7044 10906
rect 7044 10854 7090 10906
rect 6794 10852 6850 10854
rect 6874 10852 6930 10854
rect 6954 10852 7010 10854
rect 7034 10852 7090 10854
rect 7746 10648 7802 10704
rect 1852 10362 1908 10364
rect 1932 10362 1988 10364
rect 2012 10362 2068 10364
rect 2092 10362 2148 10364
rect 1852 10310 1898 10362
rect 1898 10310 1908 10362
rect 1932 10310 1962 10362
rect 1962 10310 1974 10362
rect 1974 10310 1988 10362
rect 2012 10310 2026 10362
rect 2026 10310 2038 10362
rect 2038 10310 2068 10362
rect 2092 10310 2102 10362
rect 2102 10310 2148 10362
rect 1852 10308 1908 10310
rect 1932 10308 1988 10310
rect 2012 10308 2068 10310
rect 2092 10308 2148 10310
rect 3829 10362 3885 10364
rect 3909 10362 3965 10364
rect 3989 10362 4045 10364
rect 4069 10362 4125 10364
rect 3829 10310 3875 10362
rect 3875 10310 3885 10362
rect 3909 10310 3939 10362
rect 3939 10310 3951 10362
rect 3951 10310 3965 10362
rect 3989 10310 4003 10362
rect 4003 10310 4015 10362
rect 4015 10310 4045 10362
rect 4069 10310 4079 10362
rect 4079 10310 4125 10362
rect 3829 10308 3885 10310
rect 3909 10308 3965 10310
rect 3989 10308 4045 10310
rect 4069 10308 4125 10310
rect 5806 10362 5862 10364
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 5806 10310 5852 10362
rect 5852 10310 5862 10362
rect 5886 10310 5916 10362
rect 5916 10310 5928 10362
rect 5928 10310 5942 10362
rect 5966 10310 5980 10362
rect 5980 10310 5992 10362
rect 5992 10310 6022 10362
rect 6046 10310 6056 10362
rect 6056 10310 6102 10362
rect 5806 10308 5862 10310
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 7783 10362 7839 10364
rect 7863 10362 7919 10364
rect 7943 10362 7999 10364
rect 8023 10362 8079 10364
rect 7783 10310 7829 10362
rect 7829 10310 7839 10362
rect 7863 10310 7893 10362
rect 7893 10310 7905 10362
rect 7905 10310 7919 10362
rect 7943 10310 7957 10362
rect 7957 10310 7969 10362
rect 7969 10310 7999 10362
rect 8023 10310 8033 10362
rect 8033 10310 8079 10362
rect 7783 10308 7839 10310
rect 7863 10308 7919 10310
rect 7943 10308 7999 10310
rect 8023 10308 8079 10310
rect 2840 9818 2896 9820
rect 2920 9818 2976 9820
rect 3000 9818 3056 9820
rect 3080 9818 3136 9820
rect 2840 9766 2886 9818
rect 2886 9766 2896 9818
rect 2920 9766 2950 9818
rect 2950 9766 2962 9818
rect 2962 9766 2976 9818
rect 3000 9766 3014 9818
rect 3014 9766 3026 9818
rect 3026 9766 3056 9818
rect 3080 9766 3090 9818
rect 3090 9766 3136 9818
rect 2840 9764 2896 9766
rect 2920 9764 2976 9766
rect 3000 9764 3056 9766
rect 3080 9764 3136 9766
rect 4817 9818 4873 9820
rect 4897 9818 4953 9820
rect 4977 9818 5033 9820
rect 5057 9818 5113 9820
rect 4817 9766 4863 9818
rect 4863 9766 4873 9818
rect 4897 9766 4927 9818
rect 4927 9766 4939 9818
rect 4939 9766 4953 9818
rect 4977 9766 4991 9818
rect 4991 9766 5003 9818
rect 5003 9766 5033 9818
rect 5057 9766 5067 9818
rect 5067 9766 5113 9818
rect 4817 9764 4873 9766
rect 4897 9764 4953 9766
rect 4977 9764 5033 9766
rect 5057 9764 5113 9766
rect 6794 9818 6850 9820
rect 6874 9818 6930 9820
rect 6954 9818 7010 9820
rect 7034 9818 7090 9820
rect 6794 9766 6840 9818
rect 6840 9766 6850 9818
rect 6874 9766 6904 9818
rect 6904 9766 6916 9818
rect 6916 9766 6930 9818
rect 6954 9766 6968 9818
rect 6968 9766 6980 9818
rect 6980 9766 7010 9818
rect 7034 9766 7044 9818
rect 7044 9766 7090 9818
rect 6794 9764 6850 9766
rect 6874 9764 6930 9766
rect 6954 9764 7010 9766
rect 7034 9764 7090 9766
rect 1852 9274 1908 9276
rect 1932 9274 1988 9276
rect 2012 9274 2068 9276
rect 2092 9274 2148 9276
rect 1852 9222 1898 9274
rect 1898 9222 1908 9274
rect 1932 9222 1962 9274
rect 1962 9222 1974 9274
rect 1974 9222 1988 9274
rect 2012 9222 2026 9274
rect 2026 9222 2038 9274
rect 2038 9222 2068 9274
rect 2092 9222 2102 9274
rect 2102 9222 2148 9274
rect 1852 9220 1908 9222
rect 1932 9220 1988 9222
rect 2012 9220 2068 9222
rect 2092 9220 2148 9222
rect 3829 9274 3885 9276
rect 3909 9274 3965 9276
rect 3989 9274 4045 9276
rect 4069 9274 4125 9276
rect 3829 9222 3875 9274
rect 3875 9222 3885 9274
rect 3909 9222 3939 9274
rect 3939 9222 3951 9274
rect 3951 9222 3965 9274
rect 3989 9222 4003 9274
rect 4003 9222 4015 9274
rect 4015 9222 4045 9274
rect 4069 9222 4079 9274
rect 4079 9222 4125 9274
rect 3829 9220 3885 9222
rect 3909 9220 3965 9222
rect 3989 9220 4045 9222
rect 4069 9220 4125 9222
rect 5806 9274 5862 9276
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 5806 9222 5852 9274
rect 5852 9222 5862 9274
rect 5886 9222 5916 9274
rect 5916 9222 5928 9274
rect 5928 9222 5942 9274
rect 5966 9222 5980 9274
rect 5980 9222 5992 9274
rect 5992 9222 6022 9274
rect 6046 9222 6056 9274
rect 6056 9222 6102 9274
rect 5806 9220 5862 9222
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 7783 9274 7839 9276
rect 7863 9274 7919 9276
rect 7943 9274 7999 9276
rect 8023 9274 8079 9276
rect 7783 9222 7829 9274
rect 7829 9222 7839 9274
rect 7863 9222 7893 9274
rect 7893 9222 7905 9274
rect 7905 9222 7919 9274
rect 7943 9222 7957 9274
rect 7957 9222 7969 9274
rect 7969 9222 7999 9274
rect 8023 9222 8033 9274
rect 8033 9222 8079 9274
rect 7783 9220 7839 9222
rect 7863 9220 7919 9222
rect 7943 9220 7999 9222
rect 8023 9220 8079 9222
rect 8771 10906 8827 10908
rect 8851 10906 8907 10908
rect 8931 10906 8987 10908
rect 9011 10906 9067 10908
rect 8771 10854 8817 10906
rect 8817 10854 8827 10906
rect 8851 10854 8881 10906
rect 8881 10854 8893 10906
rect 8893 10854 8907 10906
rect 8931 10854 8945 10906
rect 8945 10854 8957 10906
rect 8957 10854 8987 10906
rect 9011 10854 9021 10906
rect 9021 10854 9067 10906
rect 8771 10852 8827 10854
rect 8851 10852 8907 10854
rect 8931 10852 8987 10854
rect 9011 10852 9067 10854
rect 7838 8880 7894 8936
rect 2840 8730 2896 8732
rect 2920 8730 2976 8732
rect 3000 8730 3056 8732
rect 3080 8730 3136 8732
rect 2840 8678 2886 8730
rect 2886 8678 2896 8730
rect 2920 8678 2950 8730
rect 2950 8678 2962 8730
rect 2962 8678 2976 8730
rect 3000 8678 3014 8730
rect 3014 8678 3026 8730
rect 3026 8678 3056 8730
rect 3080 8678 3090 8730
rect 3090 8678 3136 8730
rect 2840 8676 2896 8678
rect 2920 8676 2976 8678
rect 3000 8676 3056 8678
rect 3080 8676 3136 8678
rect 4817 8730 4873 8732
rect 4897 8730 4953 8732
rect 4977 8730 5033 8732
rect 5057 8730 5113 8732
rect 4817 8678 4863 8730
rect 4863 8678 4873 8730
rect 4897 8678 4927 8730
rect 4927 8678 4939 8730
rect 4939 8678 4953 8730
rect 4977 8678 4991 8730
rect 4991 8678 5003 8730
rect 5003 8678 5033 8730
rect 5057 8678 5067 8730
rect 5067 8678 5113 8730
rect 4817 8676 4873 8678
rect 4897 8676 4953 8678
rect 4977 8676 5033 8678
rect 5057 8676 5113 8678
rect 6794 8730 6850 8732
rect 6874 8730 6930 8732
rect 6954 8730 7010 8732
rect 7034 8730 7090 8732
rect 6794 8678 6840 8730
rect 6840 8678 6850 8730
rect 6874 8678 6904 8730
rect 6904 8678 6916 8730
rect 6916 8678 6930 8730
rect 6954 8678 6968 8730
rect 6968 8678 6980 8730
rect 6980 8678 7010 8730
rect 7034 8678 7044 8730
rect 7044 8678 7090 8730
rect 6794 8676 6850 8678
rect 6874 8676 6930 8678
rect 6954 8676 7010 8678
rect 7034 8676 7090 8678
rect 1852 8186 1908 8188
rect 1932 8186 1988 8188
rect 2012 8186 2068 8188
rect 2092 8186 2148 8188
rect 1852 8134 1898 8186
rect 1898 8134 1908 8186
rect 1932 8134 1962 8186
rect 1962 8134 1974 8186
rect 1974 8134 1988 8186
rect 2012 8134 2026 8186
rect 2026 8134 2038 8186
rect 2038 8134 2068 8186
rect 2092 8134 2102 8186
rect 2102 8134 2148 8186
rect 1852 8132 1908 8134
rect 1932 8132 1988 8134
rect 2012 8132 2068 8134
rect 2092 8132 2148 8134
rect 3829 8186 3885 8188
rect 3909 8186 3965 8188
rect 3989 8186 4045 8188
rect 4069 8186 4125 8188
rect 3829 8134 3875 8186
rect 3875 8134 3885 8186
rect 3909 8134 3939 8186
rect 3939 8134 3951 8186
rect 3951 8134 3965 8186
rect 3989 8134 4003 8186
rect 4003 8134 4015 8186
rect 4015 8134 4045 8186
rect 4069 8134 4079 8186
rect 4079 8134 4125 8186
rect 3829 8132 3885 8134
rect 3909 8132 3965 8134
rect 3989 8132 4045 8134
rect 4069 8132 4125 8134
rect 5806 8186 5862 8188
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 5806 8134 5852 8186
rect 5852 8134 5862 8186
rect 5886 8134 5916 8186
rect 5916 8134 5928 8186
rect 5928 8134 5942 8186
rect 5966 8134 5980 8186
rect 5980 8134 5992 8186
rect 5992 8134 6022 8186
rect 6046 8134 6056 8186
rect 6056 8134 6102 8186
rect 5806 8132 5862 8134
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 7783 8186 7839 8188
rect 7863 8186 7919 8188
rect 7943 8186 7999 8188
rect 8023 8186 8079 8188
rect 7783 8134 7829 8186
rect 7829 8134 7839 8186
rect 7863 8134 7893 8186
rect 7893 8134 7905 8186
rect 7905 8134 7919 8186
rect 7943 8134 7957 8186
rect 7957 8134 7969 8186
rect 7969 8134 7999 8186
rect 8023 8134 8033 8186
rect 8033 8134 8079 8186
rect 7783 8132 7839 8134
rect 7863 8132 7919 8134
rect 7943 8132 7999 8134
rect 8023 8132 8079 8134
rect 2840 7642 2896 7644
rect 2920 7642 2976 7644
rect 3000 7642 3056 7644
rect 3080 7642 3136 7644
rect 2840 7590 2886 7642
rect 2886 7590 2896 7642
rect 2920 7590 2950 7642
rect 2950 7590 2962 7642
rect 2962 7590 2976 7642
rect 3000 7590 3014 7642
rect 3014 7590 3026 7642
rect 3026 7590 3056 7642
rect 3080 7590 3090 7642
rect 3090 7590 3136 7642
rect 2840 7588 2896 7590
rect 2920 7588 2976 7590
rect 3000 7588 3056 7590
rect 3080 7588 3136 7590
rect 4817 7642 4873 7644
rect 4897 7642 4953 7644
rect 4977 7642 5033 7644
rect 5057 7642 5113 7644
rect 4817 7590 4863 7642
rect 4863 7590 4873 7642
rect 4897 7590 4927 7642
rect 4927 7590 4939 7642
rect 4939 7590 4953 7642
rect 4977 7590 4991 7642
rect 4991 7590 5003 7642
rect 5003 7590 5033 7642
rect 5057 7590 5067 7642
rect 5067 7590 5113 7642
rect 4817 7588 4873 7590
rect 4897 7588 4953 7590
rect 4977 7588 5033 7590
rect 5057 7588 5113 7590
rect 6794 7642 6850 7644
rect 6874 7642 6930 7644
rect 6954 7642 7010 7644
rect 7034 7642 7090 7644
rect 6794 7590 6840 7642
rect 6840 7590 6850 7642
rect 6874 7590 6904 7642
rect 6904 7590 6916 7642
rect 6916 7590 6930 7642
rect 6954 7590 6968 7642
rect 6968 7590 6980 7642
rect 6980 7590 7010 7642
rect 7034 7590 7044 7642
rect 7044 7590 7090 7642
rect 6794 7588 6850 7590
rect 6874 7588 6930 7590
rect 6954 7588 7010 7590
rect 7034 7588 7090 7590
rect 1852 7098 1908 7100
rect 1932 7098 1988 7100
rect 2012 7098 2068 7100
rect 2092 7098 2148 7100
rect 1852 7046 1898 7098
rect 1898 7046 1908 7098
rect 1932 7046 1962 7098
rect 1962 7046 1974 7098
rect 1974 7046 1988 7098
rect 2012 7046 2026 7098
rect 2026 7046 2038 7098
rect 2038 7046 2068 7098
rect 2092 7046 2102 7098
rect 2102 7046 2148 7098
rect 1852 7044 1908 7046
rect 1932 7044 1988 7046
rect 2012 7044 2068 7046
rect 2092 7044 2148 7046
rect 3829 7098 3885 7100
rect 3909 7098 3965 7100
rect 3989 7098 4045 7100
rect 4069 7098 4125 7100
rect 3829 7046 3875 7098
rect 3875 7046 3885 7098
rect 3909 7046 3939 7098
rect 3939 7046 3951 7098
rect 3951 7046 3965 7098
rect 3989 7046 4003 7098
rect 4003 7046 4015 7098
rect 4015 7046 4045 7098
rect 4069 7046 4079 7098
rect 4079 7046 4125 7098
rect 3829 7044 3885 7046
rect 3909 7044 3965 7046
rect 3989 7044 4045 7046
rect 4069 7044 4125 7046
rect 5806 7098 5862 7100
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 5806 7046 5852 7098
rect 5852 7046 5862 7098
rect 5886 7046 5916 7098
rect 5916 7046 5928 7098
rect 5928 7046 5942 7098
rect 5966 7046 5980 7098
rect 5980 7046 5992 7098
rect 5992 7046 6022 7098
rect 6046 7046 6056 7098
rect 6056 7046 6102 7098
rect 5806 7044 5862 7046
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 7783 7098 7839 7100
rect 7863 7098 7919 7100
rect 7943 7098 7999 7100
rect 8023 7098 8079 7100
rect 7783 7046 7829 7098
rect 7829 7046 7839 7098
rect 7863 7046 7893 7098
rect 7893 7046 7905 7098
rect 7905 7046 7919 7098
rect 7943 7046 7957 7098
rect 7957 7046 7969 7098
rect 7969 7046 7999 7098
rect 8023 7046 8033 7098
rect 8033 7046 8079 7098
rect 7783 7044 7839 7046
rect 7863 7044 7919 7046
rect 7943 7044 7999 7046
rect 8023 7044 8079 7046
rect 7838 6840 7894 6896
rect 8771 9818 8827 9820
rect 8851 9818 8907 9820
rect 8931 9818 8987 9820
rect 9011 9818 9067 9820
rect 8771 9766 8817 9818
rect 8817 9766 8827 9818
rect 8851 9766 8881 9818
rect 8881 9766 8893 9818
rect 8893 9766 8907 9818
rect 8931 9766 8945 9818
rect 8945 9766 8957 9818
rect 8957 9766 8987 9818
rect 9011 9766 9021 9818
rect 9021 9766 9067 9818
rect 8771 9764 8827 9766
rect 8851 9764 8907 9766
rect 8931 9764 8987 9766
rect 9011 9764 9067 9766
rect 8771 8730 8827 8732
rect 8851 8730 8907 8732
rect 8931 8730 8987 8732
rect 9011 8730 9067 8732
rect 8771 8678 8817 8730
rect 8817 8678 8827 8730
rect 8851 8678 8881 8730
rect 8881 8678 8893 8730
rect 8893 8678 8907 8730
rect 8931 8678 8945 8730
rect 8945 8678 8957 8730
rect 8957 8678 8987 8730
rect 9011 8678 9021 8730
rect 9021 8678 9067 8730
rect 8771 8676 8827 8678
rect 8851 8676 8907 8678
rect 8931 8676 8987 8678
rect 9011 8676 9067 8678
rect 8771 7642 8827 7644
rect 8851 7642 8907 7644
rect 8931 7642 8987 7644
rect 9011 7642 9067 7644
rect 8771 7590 8817 7642
rect 8817 7590 8827 7642
rect 8851 7590 8881 7642
rect 8881 7590 8893 7642
rect 8893 7590 8907 7642
rect 8931 7590 8945 7642
rect 8945 7590 8957 7642
rect 8957 7590 8987 7642
rect 9011 7590 9021 7642
rect 9021 7590 9067 7642
rect 8771 7588 8827 7590
rect 8851 7588 8907 7590
rect 8931 7588 8987 7590
rect 9011 7588 9067 7590
rect 2840 6554 2896 6556
rect 2920 6554 2976 6556
rect 3000 6554 3056 6556
rect 3080 6554 3136 6556
rect 2840 6502 2886 6554
rect 2886 6502 2896 6554
rect 2920 6502 2950 6554
rect 2950 6502 2962 6554
rect 2962 6502 2976 6554
rect 3000 6502 3014 6554
rect 3014 6502 3026 6554
rect 3026 6502 3056 6554
rect 3080 6502 3090 6554
rect 3090 6502 3136 6554
rect 2840 6500 2896 6502
rect 2920 6500 2976 6502
rect 3000 6500 3056 6502
rect 3080 6500 3136 6502
rect 4817 6554 4873 6556
rect 4897 6554 4953 6556
rect 4977 6554 5033 6556
rect 5057 6554 5113 6556
rect 4817 6502 4863 6554
rect 4863 6502 4873 6554
rect 4897 6502 4927 6554
rect 4927 6502 4939 6554
rect 4939 6502 4953 6554
rect 4977 6502 4991 6554
rect 4991 6502 5003 6554
rect 5003 6502 5033 6554
rect 5057 6502 5067 6554
rect 5067 6502 5113 6554
rect 4817 6500 4873 6502
rect 4897 6500 4953 6502
rect 4977 6500 5033 6502
rect 5057 6500 5113 6502
rect 6794 6554 6850 6556
rect 6874 6554 6930 6556
rect 6954 6554 7010 6556
rect 7034 6554 7090 6556
rect 6794 6502 6840 6554
rect 6840 6502 6850 6554
rect 6874 6502 6904 6554
rect 6904 6502 6916 6554
rect 6916 6502 6930 6554
rect 6954 6502 6968 6554
rect 6968 6502 6980 6554
rect 6980 6502 7010 6554
rect 7034 6502 7044 6554
rect 7044 6502 7090 6554
rect 6794 6500 6850 6502
rect 6874 6500 6930 6502
rect 6954 6500 7010 6502
rect 7034 6500 7090 6502
rect 1852 6010 1908 6012
rect 1932 6010 1988 6012
rect 2012 6010 2068 6012
rect 2092 6010 2148 6012
rect 1852 5958 1898 6010
rect 1898 5958 1908 6010
rect 1932 5958 1962 6010
rect 1962 5958 1974 6010
rect 1974 5958 1988 6010
rect 2012 5958 2026 6010
rect 2026 5958 2038 6010
rect 2038 5958 2068 6010
rect 2092 5958 2102 6010
rect 2102 5958 2148 6010
rect 1852 5956 1908 5958
rect 1932 5956 1988 5958
rect 2012 5956 2068 5958
rect 2092 5956 2148 5958
rect 3829 6010 3885 6012
rect 3909 6010 3965 6012
rect 3989 6010 4045 6012
rect 4069 6010 4125 6012
rect 3829 5958 3875 6010
rect 3875 5958 3885 6010
rect 3909 5958 3939 6010
rect 3939 5958 3951 6010
rect 3951 5958 3965 6010
rect 3989 5958 4003 6010
rect 4003 5958 4015 6010
rect 4015 5958 4045 6010
rect 4069 5958 4079 6010
rect 4079 5958 4125 6010
rect 3829 5956 3885 5958
rect 3909 5956 3965 5958
rect 3989 5956 4045 5958
rect 4069 5956 4125 5958
rect 5806 6010 5862 6012
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 5806 5958 5852 6010
rect 5852 5958 5862 6010
rect 5886 5958 5916 6010
rect 5916 5958 5928 6010
rect 5928 5958 5942 6010
rect 5966 5958 5980 6010
rect 5980 5958 5992 6010
rect 5992 5958 6022 6010
rect 6046 5958 6056 6010
rect 6056 5958 6102 6010
rect 5806 5956 5862 5958
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 7783 6010 7839 6012
rect 7863 6010 7919 6012
rect 7943 6010 7999 6012
rect 8023 6010 8079 6012
rect 7783 5958 7829 6010
rect 7829 5958 7839 6010
rect 7863 5958 7893 6010
rect 7893 5958 7905 6010
rect 7905 5958 7919 6010
rect 7943 5958 7957 6010
rect 7957 5958 7969 6010
rect 7969 5958 7999 6010
rect 8023 5958 8033 6010
rect 8033 5958 8079 6010
rect 7783 5956 7839 5958
rect 7863 5956 7919 5958
rect 7943 5956 7999 5958
rect 8023 5956 8079 5958
rect 2840 5466 2896 5468
rect 2920 5466 2976 5468
rect 3000 5466 3056 5468
rect 3080 5466 3136 5468
rect 2840 5414 2886 5466
rect 2886 5414 2896 5466
rect 2920 5414 2950 5466
rect 2950 5414 2962 5466
rect 2962 5414 2976 5466
rect 3000 5414 3014 5466
rect 3014 5414 3026 5466
rect 3026 5414 3056 5466
rect 3080 5414 3090 5466
rect 3090 5414 3136 5466
rect 2840 5412 2896 5414
rect 2920 5412 2976 5414
rect 3000 5412 3056 5414
rect 3080 5412 3136 5414
rect 4817 5466 4873 5468
rect 4897 5466 4953 5468
rect 4977 5466 5033 5468
rect 5057 5466 5113 5468
rect 4817 5414 4863 5466
rect 4863 5414 4873 5466
rect 4897 5414 4927 5466
rect 4927 5414 4939 5466
rect 4939 5414 4953 5466
rect 4977 5414 4991 5466
rect 4991 5414 5003 5466
rect 5003 5414 5033 5466
rect 5057 5414 5067 5466
rect 5067 5414 5113 5466
rect 4817 5412 4873 5414
rect 4897 5412 4953 5414
rect 4977 5412 5033 5414
rect 5057 5412 5113 5414
rect 6794 5466 6850 5468
rect 6874 5466 6930 5468
rect 6954 5466 7010 5468
rect 7034 5466 7090 5468
rect 6794 5414 6840 5466
rect 6840 5414 6850 5466
rect 6874 5414 6904 5466
rect 6904 5414 6916 5466
rect 6916 5414 6930 5466
rect 6954 5414 6968 5466
rect 6968 5414 6980 5466
rect 6980 5414 7010 5466
rect 7034 5414 7044 5466
rect 7044 5414 7090 5466
rect 6794 5412 6850 5414
rect 6874 5412 6930 5414
rect 6954 5412 7010 5414
rect 7034 5412 7090 5414
rect 8771 6554 8827 6556
rect 8851 6554 8907 6556
rect 8931 6554 8987 6556
rect 9011 6554 9067 6556
rect 8771 6502 8817 6554
rect 8817 6502 8827 6554
rect 8851 6502 8881 6554
rect 8881 6502 8893 6554
rect 8893 6502 8907 6554
rect 8931 6502 8945 6554
rect 8945 6502 8957 6554
rect 8957 6502 8987 6554
rect 9011 6502 9021 6554
rect 9021 6502 9067 6554
rect 8771 6500 8827 6502
rect 8851 6500 8907 6502
rect 8931 6500 8987 6502
rect 9011 6500 9067 6502
rect 8771 5466 8827 5468
rect 8851 5466 8907 5468
rect 8931 5466 8987 5468
rect 9011 5466 9067 5468
rect 8771 5414 8817 5466
rect 8817 5414 8827 5466
rect 8851 5414 8881 5466
rect 8881 5414 8893 5466
rect 8893 5414 8907 5466
rect 8931 5414 8945 5466
rect 8945 5414 8957 5466
rect 8957 5414 8987 5466
rect 9011 5414 9021 5466
rect 9021 5414 9067 5466
rect 8771 5412 8827 5414
rect 8851 5412 8907 5414
rect 8931 5412 8987 5414
rect 9011 5412 9067 5414
rect 8206 4972 8208 4992
rect 8208 4972 8260 4992
rect 8260 4972 8262 4992
rect 8206 4936 8262 4972
rect 1852 4922 1908 4924
rect 1932 4922 1988 4924
rect 2012 4922 2068 4924
rect 2092 4922 2148 4924
rect 1852 4870 1898 4922
rect 1898 4870 1908 4922
rect 1932 4870 1962 4922
rect 1962 4870 1974 4922
rect 1974 4870 1988 4922
rect 2012 4870 2026 4922
rect 2026 4870 2038 4922
rect 2038 4870 2068 4922
rect 2092 4870 2102 4922
rect 2102 4870 2148 4922
rect 1852 4868 1908 4870
rect 1932 4868 1988 4870
rect 2012 4868 2068 4870
rect 2092 4868 2148 4870
rect 3829 4922 3885 4924
rect 3909 4922 3965 4924
rect 3989 4922 4045 4924
rect 4069 4922 4125 4924
rect 3829 4870 3875 4922
rect 3875 4870 3885 4922
rect 3909 4870 3939 4922
rect 3939 4870 3951 4922
rect 3951 4870 3965 4922
rect 3989 4870 4003 4922
rect 4003 4870 4015 4922
rect 4015 4870 4045 4922
rect 4069 4870 4079 4922
rect 4079 4870 4125 4922
rect 3829 4868 3885 4870
rect 3909 4868 3965 4870
rect 3989 4868 4045 4870
rect 4069 4868 4125 4870
rect 5806 4922 5862 4924
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 5806 4870 5852 4922
rect 5852 4870 5862 4922
rect 5886 4870 5916 4922
rect 5916 4870 5928 4922
rect 5928 4870 5942 4922
rect 5966 4870 5980 4922
rect 5980 4870 5992 4922
rect 5992 4870 6022 4922
rect 6046 4870 6056 4922
rect 6056 4870 6102 4922
rect 5806 4868 5862 4870
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 7783 4922 7839 4924
rect 7863 4922 7919 4924
rect 7943 4922 7999 4924
rect 8023 4922 8079 4924
rect 7783 4870 7829 4922
rect 7829 4870 7839 4922
rect 7863 4870 7893 4922
rect 7893 4870 7905 4922
rect 7905 4870 7919 4922
rect 7943 4870 7957 4922
rect 7957 4870 7969 4922
rect 7969 4870 7999 4922
rect 8023 4870 8033 4922
rect 8033 4870 8079 4922
rect 7783 4868 7839 4870
rect 7863 4868 7919 4870
rect 7943 4868 7999 4870
rect 8023 4868 8079 4870
rect 2840 4378 2896 4380
rect 2920 4378 2976 4380
rect 3000 4378 3056 4380
rect 3080 4378 3136 4380
rect 2840 4326 2886 4378
rect 2886 4326 2896 4378
rect 2920 4326 2950 4378
rect 2950 4326 2962 4378
rect 2962 4326 2976 4378
rect 3000 4326 3014 4378
rect 3014 4326 3026 4378
rect 3026 4326 3056 4378
rect 3080 4326 3090 4378
rect 3090 4326 3136 4378
rect 2840 4324 2896 4326
rect 2920 4324 2976 4326
rect 3000 4324 3056 4326
rect 3080 4324 3136 4326
rect 4817 4378 4873 4380
rect 4897 4378 4953 4380
rect 4977 4378 5033 4380
rect 5057 4378 5113 4380
rect 4817 4326 4863 4378
rect 4863 4326 4873 4378
rect 4897 4326 4927 4378
rect 4927 4326 4939 4378
rect 4939 4326 4953 4378
rect 4977 4326 4991 4378
rect 4991 4326 5003 4378
rect 5003 4326 5033 4378
rect 5057 4326 5067 4378
rect 5067 4326 5113 4378
rect 4817 4324 4873 4326
rect 4897 4324 4953 4326
rect 4977 4324 5033 4326
rect 5057 4324 5113 4326
rect 6794 4378 6850 4380
rect 6874 4378 6930 4380
rect 6954 4378 7010 4380
rect 7034 4378 7090 4380
rect 6794 4326 6840 4378
rect 6840 4326 6850 4378
rect 6874 4326 6904 4378
rect 6904 4326 6916 4378
rect 6916 4326 6930 4378
rect 6954 4326 6968 4378
rect 6968 4326 6980 4378
rect 6980 4326 7010 4378
rect 7034 4326 7044 4378
rect 7044 4326 7090 4378
rect 6794 4324 6850 4326
rect 6874 4324 6930 4326
rect 6954 4324 7010 4326
rect 7034 4324 7090 4326
rect 1852 3834 1908 3836
rect 1932 3834 1988 3836
rect 2012 3834 2068 3836
rect 2092 3834 2148 3836
rect 1852 3782 1898 3834
rect 1898 3782 1908 3834
rect 1932 3782 1962 3834
rect 1962 3782 1974 3834
rect 1974 3782 1988 3834
rect 2012 3782 2026 3834
rect 2026 3782 2038 3834
rect 2038 3782 2068 3834
rect 2092 3782 2102 3834
rect 2102 3782 2148 3834
rect 1852 3780 1908 3782
rect 1932 3780 1988 3782
rect 2012 3780 2068 3782
rect 2092 3780 2148 3782
rect 3829 3834 3885 3836
rect 3909 3834 3965 3836
rect 3989 3834 4045 3836
rect 4069 3834 4125 3836
rect 3829 3782 3875 3834
rect 3875 3782 3885 3834
rect 3909 3782 3939 3834
rect 3939 3782 3951 3834
rect 3951 3782 3965 3834
rect 3989 3782 4003 3834
rect 4003 3782 4015 3834
rect 4015 3782 4045 3834
rect 4069 3782 4079 3834
rect 4079 3782 4125 3834
rect 3829 3780 3885 3782
rect 3909 3780 3965 3782
rect 3989 3780 4045 3782
rect 4069 3780 4125 3782
rect 5806 3834 5862 3836
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 5806 3782 5852 3834
rect 5852 3782 5862 3834
rect 5886 3782 5916 3834
rect 5916 3782 5928 3834
rect 5928 3782 5942 3834
rect 5966 3782 5980 3834
rect 5980 3782 5992 3834
rect 5992 3782 6022 3834
rect 6046 3782 6056 3834
rect 6056 3782 6102 3834
rect 5806 3780 5862 3782
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 7783 3834 7839 3836
rect 7863 3834 7919 3836
rect 7943 3834 7999 3836
rect 8023 3834 8079 3836
rect 7783 3782 7829 3834
rect 7829 3782 7839 3834
rect 7863 3782 7893 3834
rect 7893 3782 7905 3834
rect 7905 3782 7919 3834
rect 7943 3782 7957 3834
rect 7957 3782 7969 3834
rect 7969 3782 7999 3834
rect 8023 3782 8033 3834
rect 8033 3782 8079 3834
rect 7783 3780 7839 3782
rect 7863 3780 7919 3782
rect 7943 3780 7999 3782
rect 8023 3780 8079 3782
rect 2840 3290 2896 3292
rect 2920 3290 2976 3292
rect 3000 3290 3056 3292
rect 3080 3290 3136 3292
rect 2840 3238 2886 3290
rect 2886 3238 2896 3290
rect 2920 3238 2950 3290
rect 2950 3238 2962 3290
rect 2962 3238 2976 3290
rect 3000 3238 3014 3290
rect 3014 3238 3026 3290
rect 3026 3238 3056 3290
rect 3080 3238 3090 3290
rect 3090 3238 3136 3290
rect 2840 3236 2896 3238
rect 2920 3236 2976 3238
rect 3000 3236 3056 3238
rect 3080 3236 3136 3238
rect 4817 3290 4873 3292
rect 4897 3290 4953 3292
rect 4977 3290 5033 3292
rect 5057 3290 5113 3292
rect 4817 3238 4863 3290
rect 4863 3238 4873 3290
rect 4897 3238 4927 3290
rect 4927 3238 4939 3290
rect 4939 3238 4953 3290
rect 4977 3238 4991 3290
rect 4991 3238 5003 3290
rect 5003 3238 5033 3290
rect 5057 3238 5067 3290
rect 5067 3238 5113 3290
rect 4817 3236 4873 3238
rect 4897 3236 4953 3238
rect 4977 3236 5033 3238
rect 5057 3236 5113 3238
rect 6794 3290 6850 3292
rect 6874 3290 6930 3292
rect 6954 3290 7010 3292
rect 7034 3290 7090 3292
rect 6794 3238 6840 3290
rect 6840 3238 6850 3290
rect 6874 3238 6904 3290
rect 6904 3238 6916 3290
rect 6916 3238 6930 3290
rect 6954 3238 6968 3290
rect 6968 3238 6980 3290
rect 6980 3238 7010 3290
rect 7034 3238 7044 3290
rect 7044 3238 7090 3290
rect 6794 3236 6850 3238
rect 6874 3236 6930 3238
rect 6954 3236 7010 3238
rect 7034 3236 7090 3238
rect 7654 3032 7710 3088
rect 8771 4378 8827 4380
rect 8851 4378 8907 4380
rect 8931 4378 8987 4380
rect 9011 4378 9067 4380
rect 8771 4326 8817 4378
rect 8817 4326 8827 4378
rect 8851 4326 8881 4378
rect 8881 4326 8893 4378
rect 8893 4326 8907 4378
rect 8931 4326 8945 4378
rect 8945 4326 8957 4378
rect 8957 4326 8987 4378
rect 9011 4326 9021 4378
rect 9021 4326 9067 4378
rect 8771 4324 8827 4326
rect 8851 4324 8907 4326
rect 8931 4324 8987 4326
rect 9011 4324 9067 4326
rect 8771 3290 8827 3292
rect 8851 3290 8907 3292
rect 8931 3290 8987 3292
rect 9011 3290 9067 3292
rect 8771 3238 8817 3290
rect 8817 3238 8827 3290
rect 8851 3238 8881 3290
rect 8881 3238 8893 3290
rect 8893 3238 8907 3290
rect 8931 3238 8945 3290
rect 8945 3238 8957 3290
rect 8957 3238 8987 3290
rect 9011 3238 9021 3290
rect 9021 3238 9067 3290
rect 8771 3236 8827 3238
rect 8851 3236 8907 3238
rect 8931 3236 8987 3238
rect 9011 3236 9067 3238
rect 1852 2746 1908 2748
rect 1932 2746 1988 2748
rect 2012 2746 2068 2748
rect 2092 2746 2148 2748
rect 1852 2694 1898 2746
rect 1898 2694 1908 2746
rect 1932 2694 1962 2746
rect 1962 2694 1974 2746
rect 1974 2694 1988 2746
rect 2012 2694 2026 2746
rect 2026 2694 2038 2746
rect 2038 2694 2068 2746
rect 2092 2694 2102 2746
rect 2102 2694 2148 2746
rect 1852 2692 1908 2694
rect 1932 2692 1988 2694
rect 2012 2692 2068 2694
rect 2092 2692 2148 2694
rect 3829 2746 3885 2748
rect 3909 2746 3965 2748
rect 3989 2746 4045 2748
rect 4069 2746 4125 2748
rect 3829 2694 3875 2746
rect 3875 2694 3885 2746
rect 3909 2694 3939 2746
rect 3939 2694 3951 2746
rect 3951 2694 3965 2746
rect 3989 2694 4003 2746
rect 4003 2694 4015 2746
rect 4015 2694 4045 2746
rect 4069 2694 4079 2746
rect 4079 2694 4125 2746
rect 3829 2692 3885 2694
rect 3909 2692 3965 2694
rect 3989 2692 4045 2694
rect 4069 2692 4125 2694
rect 5806 2746 5862 2748
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 5806 2694 5852 2746
rect 5852 2694 5862 2746
rect 5886 2694 5916 2746
rect 5916 2694 5928 2746
rect 5928 2694 5942 2746
rect 5966 2694 5980 2746
rect 5980 2694 5992 2746
rect 5992 2694 6022 2746
rect 6046 2694 6056 2746
rect 6056 2694 6102 2746
rect 5806 2692 5862 2694
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 7783 2746 7839 2748
rect 7863 2746 7919 2748
rect 7943 2746 7999 2748
rect 8023 2746 8079 2748
rect 7783 2694 7829 2746
rect 7829 2694 7839 2746
rect 7863 2694 7893 2746
rect 7893 2694 7905 2746
rect 7905 2694 7919 2746
rect 7943 2694 7957 2746
rect 7957 2694 7969 2746
rect 7969 2694 7999 2746
rect 8023 2694 8033 2746
rect 8033 2694 8079 2746
rect 7783 2692 7839 2694
rect 7863 2692 7919 2694
rect 7943 2692 7999 2694
rect 8023 2692 8079 2694
rect 2840 2202 2896 2204
rect 2920 2202 2976 2204
rect 3000 2202 3056 2204
rect 3080 2202 3136 2204
rect 2840 2150 2886 2202
rect 2886 2150 2896 2202
rect 2920 2150 2950 2202
rect 2950 2150 2962 2202
rect 2962 2150 2976 2202
rect 3000 2150 3014 2202
rect 3014 2150 3026 2202
rect 3026 2150 3056 2202
rect 3080 2150 3090 2202
rect 3090 2150 3136 2202
rect 2840 2148 2896 2150
rect 2920 2148 2976 2150
rect 3000 2148 3056 2150
rect 3080 2148 3136 2150
rect 4817 2202 4873 2204
rect 4897 2202 4953 2204
rect 4977 2202 5033 2204
rect 5057 2202 5113 2204
rect 4817 2150 4863 2202
rect 4863 2150 4873 2202
rect 4897 2150 4927 2202
rect 4927 2150 4939 2202
rect 4939 2150 4953 2202
rect 4977 2150 4991 2202
rect 4991 2150 5003 2202
rect 5003 2150 5033 2202
rect 5057 2150 5067 2202
rect 5067 2150 5113 2202
rect 4817 2148 4873 2150
rect 4897 2148 4953 2150
rect 4977 2148 5033 2150
rect 5057 2148 5113 2150
rect 6794 2202 6850 2204
rect 6874 2202 6930 2204
rect 6954 2202 7010 2204
rect 7034 2202 7090 2204
rect 6794 2150 6840 2202
rect 6840 2150 6850 2202
rect 6874 2150 6904 2202
rect 6904 2150 6916 2202
rect 6916 2150 6930 2202
rect 6954 2150 6968 2202
rect 6968 2150 6980 2202
rect 6980 2150 7010 2202
rect 7034 2150 7044 2202
rect 7044 2150 7090 2202
rect 6794 2148 6850 2150
rect 6874 2148 6930 2150
rect 6954 2148 7010 2150
rect 7034 2148 7090 2150
rect 8771 2202 8827 2204
rect 8851 2202 8907 2204
rect 8931 2202 8987 2204
rect 9011 2202 9067 2204
rect 8771 2150 8817 2202
rect 8817 2150 8827 2202
rect 8851 2150 8881 2202
rect 8881 2150 8893 2202
rect 8893 2150 8907 2202
rect 8931 2150 8945 2202
rect 8945 2150 8957 2202
rect 8957 2150 8987 2202
rect 9011 2150 9021 2202
rect 9021 2150 9067 2202
rect 8771 2148 8827 2150
rect 8851 2148 8907 2150
rect 8931 2148 8987 2150
rect 9011 2148 9067 2150
rect 1852 1658 1908 1660
rect 1932 1658 1988 1660
rect 2012 1658 2068 1660
rect 2092 1658 2148 1660
rect 1852 1606 1898 1658
rect 1898 1606 1908 1658
rect 1932 1606 1962 1658
rect 1962 1606 1974 1658
rect 1974 1606 1988 1658
rect 2012 1606 2026 1658
rect 2026 1606 2038 1658
rect 2038 1606 2068 1658
rect 2092 1606 2102 1658
rect 2102 1606 2148 1658
rect 1852 1604 1908 1606
rect 1932 1604 1988 1606
rect 2012 1604 2068 1606
rect 2092 1604 2148 1606
rect 3829 1658 3885 1660
rect 3909 1658 3965 1660
rect 3989 1658 4045 1660
rect 4069 1658 4125 1660
rect 3829 1606 3875 1658
rect 3875 1606 3885 1658
rect 3909 1606 3939 1658
rect 3939 1606 3951 1658
rect 3951 1606 3965 1658
rect 3989 1606 4003 1658
rect 4003 1606 4015 1658
rect 4015 1606 4045 1658
rect 4069 1606 4079 1658
rect 4079 1606 4125 1658
rect 3829 1604 3885 1606
rect 3909 1604 3965 1606
rect 3989 1604 4045 1606
rect 4069 1604 4125 1606
rect 5806 1658 5862 1660
rect 5886 1658 5942 1660
rect 5966 1658 6022 1660
rect 6046 1658 6102 1660
rect 5806 1606 5852 1658
rect 5852 1606 5862 1658
rect 5886 1606 5916 1658
rect 5916 1606 5928 1658
rect 5928 1606 5942 1658
rect 5966 1606 5980 1658
rect 5980 1606 5992 1658
rect 5992 1606 6022 1658
rect 6046 1606 6056 1658
rect 6056 1606 6102 1658
rect 5806 1604 5862 1606
rect 5886 1604 5942 1606
rect 5966 1604 6022 1606
rect 6046 1604 6102 1606
rect 7783 1658 7839 1660
rect 7863 1658 7919 1660
rect 7943 1658 7999 1660
rect 8023 1658 8079 1660
rect 7783 1606 7829 1658
rect 7829 1606 7839 1658
rect 7863 1606 7893 1658
rect 7893 1606 7905 1658
rect 7905 1606 7919 1658
rect 7943 1606 7957 1658
rect 7957 1606 7969 1658
rect 7969 1606 7999 1658
rect 8023 1606 8033 1658
rect 8033 1606 8079 1658
rect 7783 1604 7839 1606
rect 7863 1604 7919 1606
rect 7943 1604 7999 1606
rect 8023 1604 8079 1606
rect 2840 1114 2896 1116
rect 2920 1114 2976 1116
rect 3000 1114 3056 1116
rect 3080 1114 3136 1116
rect 2840 1062 2886 1114
rect 2886 1062 2896 1114
rect 2920 1062 2950 1114
rect 2950 1062 2962 1114
rect 2962 1062 2976 1114
rect 3000 1062 3014 1114
rect 3014 1062 3026 1114
rect 3026 1062 3056 1114
rect 3080 1062 3090 1114
rect 3090 1062 3136 1114
rect 2840 1060 2896 1062
rect 2920 1060 2976 1062
rect 3000 1060 3056 1062
rect 3080 1060 3136 1062
rect 4817 1114 4873 1116
rect 4897 1114 4953 1116
rect 4977 1114 5033 1116
rect 5057 1114 5113 1116
rect 4817 1062 4863 1114
rect 4863 1062 4873 1114
rect 4897 1062 4927 1114
rect 4927 1062 4939 1114
rect 4939 1062 4953 1114
rect 4977 1062 4991 1114
rect 4991 1062 5003 1114
rect 5003 1062 5033 1114
rect 5057 1062 5067 1114
rect 5067 1062 5113 1114
rect 4817 1060 4873 1062
rect 4897 1060 4953 1062
rect 4977 1060 5033 1062
rect 5057 1060 5113 1062
rect 6794 1114 6850 1116
rect 6874 1114 6930 1116
rect 6954 1114 7010 1116
rect 7034 1114 7090 1116
rect 6794 1062 6840 1114
rect 6840 1062 6850 1114
rect 6874 1062 6904 1114
rect 6904 1062 6916 1114
rect 6916 1062 6930 1114
rect 6954 1062 6968 1114
rect 6968 1062 6980 1114
rect 6980 1062 7010 1114
rect 7034 1062 7044 1114
rect 7044 1062 7090 1114
rect 6794 1060 6850 1062
rect 6874 1060 6930 1062
rect 6954 1060 7010 1062
rect 7034 1060 7090 1062
rect 9310 1128 9366 1184
rect 8771 1114 8827 1116
rect 8851 1114 8907 1116
rect 8931 1114 8987 1116
rect 9011 1114 9067 1116
rect 8771 1062 8817 1114
rect 8817 1062 8827 1114
rect 8851 1062 8881 1114
rect 8881 1062 8893 1114
rect 8893 1062 8907 1114
rect 8931 1062 8945 1114
rect 8945 1062 8957 1114
rect 8957 1062 8987 1114
rect 9011 1062 9021 1114
rect 9021 1062 9067 1114
rect 8771 1060 8827 1062
rect 8851 1060 8907 1062
rect 8931 1060 8987 1062
rect 9011 1060 9067 1062
<< metal3 >>
rect 1842 14720 2158 14721
rect 1842 14656 1848 14720
rect 1912 14656 1928 14720
rect 1992 14656 2008 14720
rect 2072 14656 2088 14720
rect 2152 14656 2158 14720
rect 1842 14655 2158 14656
rect 3819 14720 4135 14721
rect 3819 14656 3825 14720
rect 3889 14656 3905 14720
rect 3969 14656 3985 14720
rect 4049 14656 4065 14720
rect 4129 14656 4135 14720
rect 3819 14655 4135 14656
rect 5796 14720 6112 14721
rect 5796 14656 5802 14720
rect 5866 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6112 14720
rect 5796 14655 6112 14656
rect 7773 14720 8089 14721
rect 7773 14656 7779 14720
rect 7843 14656 7859 14720
rect 7923 14656 7939 14720
rect 8003 14656 8019 14720
rect 8083 14656 8089 14720
rect 7773 14655 8089 14656
rect 8109 14514 8175 14517
rect 9600 14514 10000 14544
rect 8109 14512 10000 14514
rect 8109 14456 8114 14512
rect 8170 14456 10000 14512
rect 8109 14454 10000 14456
rect 8109 14451 8175 14454
rect 9600 14424 10000 14454
rect 2830 14176 3146 14177
rect 2830 14112 2836 14176
rect 2900 14112 2916 14176
rect 2980 14112 2996 14176
rect 3060 14112 3076 14176
rect 3140 14112 3146 14176
rect 2830 14111 3146 14112
rect 4807 14176 5123 14177
rect 4807 14112 4813 14176
rect 4877 14112 4893 14176
rect 4957 14112 4973 14176
rect 5037 14112 5053 14176
rect 5117 14112 5123 14176
rect 4807 14111 5123 14112
rect 6784 14176 7100 14177
rect 6784 14112 6790 14176
rect 6854 14112 6870 14176
rect 6934 14112 6950 14176
rect 7014 14112 7030 14176
rect 7094 14112 7100 14176
rect 6784 14111 7100 14112
rect 8761 14176 9077 14177
rect 8761 14112 8767 14176
rect 8831 14112 8847 14176
rect 8911 14112 8927 14176
rect 8991 14112 9007 14176
rect 9071 14112 9077 14176
rect 8761 14111 9077 14112
rect 1842 13632 2158 13633
rect 1842 13568 1848 13632
rect 1912 13568 1928 13632
rect 1992 13568 2008 13632
rect 2072 13568 2088 13632
rect 2152 13568 2158 13632
rect 1842 13567 2158 13568
rect 3819 13632 4135 13633
rect 3819 13568 3825 13632
rect 3889 13568 3905 13632
rect 3969 13568 3985 13632
rect 4049 13568 4065 13632
rect 4129 13568 4135 13632
rect 3819 13567 4135 13568
rect 5796 13632 6112 13633
rect 5796 13568 5802 13632
rect 5866 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6112 13632
rect 5796 13567 6112 13568
rect 7773 13632 8089 13633
rect 7773 13568 7779 13632
rect 7843 13568 7859 13632
rect 7923 13568 7939 13632
rect 8003 13568 8019 13632
rect 8083 13568 8089 13632
rect 7773 13567 8089 13568
rect 2830 13088 3146 13089
rect 2830 13024 2836 13088
rect 2900 13024 2916 13088
rect 2980 13024 2996 13088
rect 3060 13024 3076 13088
rect 3140 13024 3146 13088
rect 2830 13023 3146 13024
rect 4807 13088 5123 13089
rect 4807 13024 4813 13088
rect 4877 13024 4893 13088
rect 4957 13024 4973 13088
rect 5037 13024 5053 13088
rect 5117 13024 5123 13088
rect 4807 13023 5123 13024
rect 6784 13088 7100 13089
rect 6784 13024 6790 13088
rect 6854 13024 6870 13088
rect 6934 13024 6950 13088
rect 7014 13024 7030 13088
rect 7094 13024 7100 13088
rect 6784 13023 7100 13024
rect 8761 13088 9077 13089
rect 8761 13024 8767 13088
rect 8831 13024 8847 13088
rect 8911 13024 8927 13088
rect 8991 13024 9007 13088
rect 9071 13024 9077 13088
rect 8761 13023 9077 13024
rect 8201 12610 8267 12613
rect 9600 12610 10000 12640
rect 8201 12608 10000 12610
rect 8201 12552 8206 12608
rect 8262 12552 10000 12608
rect 8201 12550 10000 12552
rect 8201 12547 8267 12550
rect 1842 12544 2158 12545
rect 1842 12480 1848 12544
rect 1912 12480 1928 12544
rect 1992 12480 2008 12544
rect 2072 12480 2088 12544
rect 2152 12480 2158 12544
rect 1842 12479 2158 12480
rect 3819 12544 4135 12545
rect 3819 12480 3825 12544
rect 3889 12480 3905 12544
rect 3969 12480 3985 12544
rect 4049 12480 4065 12544
rect 4129 12480 4135 12544
rect 3819 12479 4135 12480
rect 5796 12544 6112 12545
rect 5796 12480 5802 12544
rect 5866 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6112 12544
rect 5796 12479 6112 12480
rect 7773 12544 8089 12545
rect 7773 12480 7779 12544
rect 7843 12480 7859 12544
rect 7923 12480 7939 12544
rect 8003 12480 8019 12544
rect 8083 12480 8089 12544
rect 9600 12520 10000 12550
rect 7773 12479 8089 12480
rect 2830 12000 3146 12001
rect 2830 11936 2836 12000
rect 2900 11936 2916 12000
rect 2980 11936 2996 12000
rect 3060 11936 3076 12000
rect 3140 11936 3146 12000
rect 2830 11935 3146 11936
rect 4807 12000 5123 12001
rect 4807 11936 4813 12000
rect 4877 11936 4893 12000
rect 4957 11936 4973 12000
rect 5037 11936 5053 12000
rect 5117 11936 5123 12000
rect 4807 11935 5123 11936
rect 6784 12000 7100 12001
rect 6784 11936 6790 12000
rect 6854 11936 6870 12000
rect 6934 11936 6950 12000
rect 7014 11936 7030 12000
rect 7094 11936 7100 12000
rect 6784 11935 7100 11936
rect 8761 12000 9077 12001
rect 8761 11936 8767 12000
rect 8831 11936 8847 12000
rect 8911 11936 8927 12000
rect 8991 11936 9007 12000
rect 9071 11936 9077 12000
rect 8761 11935 9077 11936
rect 1842 11456 2158 11457
rect 1842 11392 1848 11456
rect 1912 11392 1928 11456
rect 1992 11392 2008 11456
rect 2072 11392 2088 11456
rect 2152 11392 2158 11456
rect 1842 11391 2158 11392
rect 3819 11456 4135 11457
rect 3819 11392 3825 11456
rect 3889 11392 3905 11456
rect 3969 11392 3985 11456
rect 4049 11392 4065 11456
rect 4129 11392 4135 11456
rect 3819 11391 4135 11392
rect 5796 11456 6112 11457
rect 5796 11392 5802 11456
rect 5866 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6112 11456
rect 5796 11391 6112 11392
rect 7773 11456 8089 11457
rect 7773 11392 7779 11456
rect 7843 11392 7859 11456
rect 7923 11392 7939 11456
rect 8003 11392 8019 11456
rect 8083 11392 8089 11456
rect 7773 11391 8089 11392
rect 2830 10912 3146 10913
rect 2830 10848 2836 10912
rect 2900 10848 2916 10912
rect 2980 10848 2996 10912
rect 3060 10848 3076 10912
rect 3140 10848 3146 10912
rect 2830 10847 3146 10848
rect 4807 10912 5123 10913
rect 4807 10848 4813 10912
rect 4877 10848 4893 10912
rect 4957 10848 4973 10912
rect 5037 10848 5053 10912
rect 5117 10848 5123 10912
rect 4807 10847 5123 10848
rect 6784 10912 7100 10913
rect 6784 10848 6790 10912
rect 6854 10848 6870 10912
rect 6934 10848 6950 10912
rect 7014 10848 7030 10912
rect 7094 10848 7100 10912
rect 6784 10847 7100 10848
rect 8761 10912 9077 10913
rect 8761 10848 8767 10912
rect 8831 10848 8847 10912
rect 8911 10848 8927 10912
rect 8991 10848 9007 10912
rect 9071 10848 9077 10912
rect 8761 10847 9077 10848
rect 7741 10706 7807 10709
rect 9600 10706 10000 10736
rect 7741 10704 10000 10706
rect 7741 10648 7746 10704
rect 7802 10648 10000 10704
rect 7741 10646 10000 10648
rect 7741 10643 7807 10646
rect 9600 10616 10000 10646
rect 1842 10368 2158 10369
rect 1842 10304 1848 10368
rect 1912 10304 1928 10368
rect 1992 10304 2008 10368
rect 2072 10304 2088 10368
rect 2152 10304 2158 10368
rect 1842 10303 2158 10304
rect 3819 10368 4135 10369
rect 3819 10304 3825 10368
rect 3889 10304 3905 10368
rect 3969 10304 3985 10368
rect 4049 10304 4065 10368
rect 4129 10304 4135 10368
rect 3819 10303 4135 10304
rect 5796 10368 6112 10369
rect 5796 10304 5802 10368
rect 5866 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6112 10368
rect 5796 10303 6112 10304
rect 7773 10368 8089 10369
rect 7773 10304 7779 10368
rect 7843 10304 7859 10368
rect 7923 10304 7939 10368
rect 8003 10304 8019 10368
rect 8083 10304 8089 10368
rect 7773 10303 8089 10304
rect 2830 9824 3146 9825
rect 2830 9760 2836 9824
rect 2900 9760 2916 9824
rect 2980 9760 2996 9824
rect 3060 9760 3076 9824
rect 3140 9760 3146 9824
rect 2830 9759 3146 9760
rect 4807 9824 5123 9825
rect 4807 9760 4813 9824
rect 4877 9760 4893 9824
rect 4957 9760 4973 9824
rect 5037 9760 5053 9824
rect 5117 9760 5123 9824
rect 4807 9759 5123 9760
rect 6784 9824 7100 9825
rect 6784 9760 6790 9824
rect 6854 9760 6870 9824
rect 6934 9760 6950 9824
rect 7014 9760 7030 9824
rect 7094 9760 7100 9824
rect 6784 9759 7100 9760
rect 8761 9824 9077 9825
rect 8761 9760 8767 9824
rect 8831 9760 8847 9824
rect 8911 9760 8927 9824
rect 8991 9760 9007 9824
rect 9071 9760 9077 9824
rect 8761 9759 9077 9760
rect 1842 9280 2158 9281
rect 1842 9216 1848 9280
rect 1912 9216 1928 9280
rect 1992 9216 2008 9280
rect 2072 9216 2088 9280
rect 2152 9216 2158 9280
rect 1842 9215 2158 9216
rect 3819 9280 4135 9281
rect 3819 9216 3825 9280
rect 3889 9216 3905 9280
rect 3969 9216 3985 9280
rect 4049 9216 4065 9280
rect 4129 9216 4135 9280
rect 3819 9215 4135 9216
rect 5796 9280 6112 9281
rect 5796 9216 5802 9280
rect 5866 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6112 9280
rect 5796 9215 6112 9216
rect 7773 9280 8089 9281
rect 7773 9216 7779 9280
rect 7843 9216 7859 9280
rect 7923 9216 7939 9280
rect 8003 9216 8019 9280
rect 8083 9216 8089 9280
rect 7773 9215 8089 9216
rect 7833 8938 7899 8941
rect 7833 8936 9322 8938
rect 7833 8880 7838 8936
rect 7894 8880 9322 8936
rect 7833 8878 9322 8880
rect 7833 8875 7899 8878
rect 9262 8802 9322 8878
rect 9600 8802 10000 8832
rect 9262 8742 10000 8802
rect 2830 8736 3146 8737
rect 2830 8672 2836 8736
rect 2900 8672 2916 8736
rect 2980 8672 2996 8736
rect 3060 8672 3076 8736
rect 3140 8672 3146 8736
rect 2830 8671 3146 8672
rect 4807 8736 5123 8737
rect 4807 8672 4813 8736
rect 4877 8672 4893 8736
rect 4957 8672 4973 8736
rect 5037 8672 5053 8736
rect 5117 8672 5123 8736
rect 4807 8671 5123 8672
rect 6784 8736 7100 8737
rect 6784 8672 6790 8736
rect 6854 8672 6870 8736
rect 6934 8672 6950 8736
rect 7014 8672 7030 8736
rect 7094 8672 7100 8736
rect 6784 8671 7100 8672
rect 8761 8736 9077 8737
rect 8761 8672 8767 8736
rect 8831 8672 8847 8736
rect 8911 8672 8927 8736
rect 8991 8672 9007 8736
rect 9071 8672 9077 8736
rect 9600 8712 10000 8742
rect 8761 8671 9077 8672
rect 1842 8192 2158 8193
rect 1842 8128 1848 8192
rect 1912 8128 1928 8192
rect 1992 8128 2008 8192
rect 2072 8128 2088 8192
rect 2152 8128 2158 8192
rect 1842 8127 2158 8128
rect 3819 8192 4135 8193
rect 3819 8128 3825 8192
rect 3889 8128 3905 8192
rect 3969 8128 3985 8192
rect 4049 8128 4065 8192
rect 4129 8128 4135 8192
rect 3819 8127 4135 8128
rect 5796 8192 6112 8193
rect 5796 8128 5802 8192
rect 5866 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6112 8192
rect 5796 8127 6112 8128
rect 7773 8192 8089 8193
rect 7773 8128 7779 8192
rect 7843 8128 7859 8192
rect 7923 8128 7939 8192
rect 8003 8128 8019 8192
rect 8083 8128 8089 8192
rect 7773 8127 8089 8128
rect 2830 7648 3146 7649
rect 2830 7584 2836 7648
rect 2900 7584 2916 7648
rect 2980 7584 2996 7648
rect 3060 7584 3076 7648
rect 3140 7584 3146 7648
rect 2830 7583 3146 7584
rect 4807 7648 5123 7649
rect 4807 7584 4813 7648
rect 4877 7584 4893 7648
rect 4957 7584 4973 7648
rect 5037 7584 5053 7648
rect 5117 7584 5123 7648
rect 4807 7583 5123 7584
rect 6784 7648 7100 7649
rect 6784 7584 6790 7648
rect 6854 7584 6870 7648
rect 6934 7584 6950 7648
rect 7014 7584 7030 7648
rect 7094 7584 7100 7648
rect 6784 7583 7100 7584
rect 8761 7648 9077 7649
rect 8761 7584 8767 7648
rect 8831 7584 8847 7648
rect 8911 7584 8927 7648
rect 8991 7584 9007 7648
rect 9071 7584 9077 7648
rect 8761 7583 9077 7584
rect 1842 7104 2158 7105
rect 1842 7040 1848 7104
rect 1912 7040 1928 7104
rect 1992 7040 2008 7104
rect 2072 7040 2088 7104
rect 2152 7040 2158 7104
rect 1842 7039 2158 7040
rect 3819 7104 4135 7105
rect 3819 7040 3825 7104
rect 3889 7040 3905 7104
rect 3969 7040 3985 7104
rect 4049 7040 4065 7104
rect 4129 7040 4135 7104
rect 3819 7039 4135 7040
rect 5796 7104 6112 7105
rect 5796 7040 5802 7104
rect 5866 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6112 7104
rect 5796 7039 6112 7040
rect 7773 7104 8089 7105
rect 7773 7040 7779 7104
rect 7843 7040 7859 7104
rect 7923 7040 7939 7104
rect 8003 7040 8019 7104
rect 8083 7040 8089 7104
rect 7773 7039 8089 7040
rect 7833 6898 7899 6901
rect 9600 6898 10000 6928
rect 7833 6896 10000 6898
rect 7833 6840 7838 6896
rect 7894 6840 10000 6896
rect 7833 6838 10000 6840
rect 7833 6835 7899 6838
rect 9600 6808 10000 6838
rect 2830 6560 3146 6561
rect 2830 6496 2836 6560
rect 2900 6496 2916 6560
rect 2980 6496 2996 6560
rect 3060 6496 3076 6560
rect 3140 6496 3146 6560
rect 2830 6495 3146 6496
rect 4807 6560 5123 6561
rect 4807 6496 4813 6560
rect 4877 6496 4893 6560
rect 4957 6496 4973 6560
rect 5037 6496 5053 6560
rect 5117 6496 5123 6560
rect 4807 6495 5123 6496
rect 6784 6560 7100 6561
rect 6784 6496 6790 6560
rect 6854 6496 6870 6560
rect 6934 6496 6950 6560
rect 7014 6496 7030 6560
rect 7094 6496 7100 6560
rect 6784 6495 7100 6496
rect 8761 6560 9077 6561
rect 8761 6496 8767 6560
rect 8831 6496 8847 6560
rect 8911 6496 8927 6560
rect 8991 6496 9007 6560
rect 9071 6496 9077 6560
rect 8761 6495 9077 6496
rect 1842 6016 2158 6017
rect 1842 5952 1848 6016
rect 1912 5952 1928 6016
rect 1992 5952 2008 6016
rect 2072 5952 2088 6016
rect 2152 5952 2158 6016
rect 1842 5951 2158 5952
rect 3819 6016 4135 6017
rect 3819 5952 3825 6016
rect 3889 5952 3905 6016
rect 3969 5952 3985 6016
rect 4049 5952 4065 6016
rect 4129 5952 4135 6016
rect 3819 5951 4135 5952
rect 5796 6016 6112 6017
rect 5796 5952 5802 6016
rect 5866 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6112 6016
rect 5796 5951 6112 5952
rect 7773 6016 8089 6017
rect 7773 5952 7779 6016
rect 7843 5952 7859 6016
rect 7923 5952 7939 6016
rect 8003 5952 8019 6016
rect 8083 5952 8089 6016
rect 7773 5951 8089 5952
rect 2830 5472 3146 5473
rect 2830 5408 2836 5472
rect 2900 5408 2916 5472
rect 2980 5408 2996 5472
rect 3060 5408 3076 5472
rect 3140 5408 3146 5472
rect 2830 5407 3146 5408
rect 4807 5472 5123 5473
rect 4807 5408 4813 5472
rect 4877 5408 4893 5472
rect 4957 5408 4973 5472
rect 5037 5408 5053 5472
rect 5117 5408 5123 5472
rect 4807 5407 5123 5408
rect 6784 5472 7100 5473
rect 6784 5408 6790 5472
rect 6854 5408 6870 5472
rect 6934 5408 6950 5472
rect 7014 5408 7030 5472
rect 7094 5408 7100 5472
rect 6784 5407 7100 5408
rect 8761 5472 9077 5473
rect 8761 5408 8767 5472
rect 8831 5408 8847 5472
rect 8911 5408 8927 5472
rect 8991 5408 9007 5472
rect 9071 5408 9077 5472
rect 8761 5407 9077 5408
rect 8201 4994 8267 4997
rect 9600 4994 10000 5024
rect 8201 4992 10000 4994
rect 8201 4936 8206 4992
rect 8262 4936 10000 4992
rect 8201 4934 10000 4936
rect 8201 4931 8267 4934
rect 1842 4928 2158 4929
rect 1842 4864 1848 4928
rect 1912 4864 1928 4928
rect 1992 4864 2008 4928
rect 2072 4864 2088 4928
rect 2152 4864 2158 4928
rect 1842 4863 2158 4864
rect 3819 4928 4135 4929
rect 3819 4864 3825 4928
rect 3889 4864 3905 4928
rect 3969 4864 3985 4928
rect 4049 4864 4065 4928
rect 4129 4864 4135 4928
rect 3819 4863 4135 4864
rect 5796 4928 6112 4929
rect 5796 4864 5802 4928
rect 5866 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6112 4928
rect 5796 4863 6112 4864
rect 7773 4928 8089 4929
rect 7773 4864 7779 4928
rect 7843 4864 7859 4928
rect 7923 4864 7939 4928
rect 8003 4864 8019 4928
rect 8083 4864 8089 4928
rect 9600 4904 10000 4934
rect 7773 4863 8089 4864
rect 2830 4384 3146 4385
rect 2830 4320 2836 4384
rect 2900 4320 2916 4384
rect 2980 4320 2996 4384
rect 3060 4320 3076 4384
rect 3140 4320 3146 4384
rect 2830 4319 3146 4320
rect 4807 4384 5123 4385
rect 4807 4320 4813 4384
rect 4877 4320 4893 4384
rect 4957 4320 4973 4384
rect 5037 4320 5053 4384
rect 5117 4320 5123 4384
rect 4807 4319 5123 4320
rect 6784 4384 7100 4385
rect 6784 4320 6790 4384
rect 6854 4320 6870 4384
rect 6934 4320 6950 4384
rect 7014 4320 7030 4384
rect 7094 4320 7100 4384
rect 6784 4319 7100 4320
rect 8761 4384 9077 4385
rect 8761 4320 8767 4384
rect 8831 4320 8847 4384
rect 8911 4320 8927 4384
rect 8991 4320 9007 4384
rect 9071 4320 9077 4384
rect 8761 4319 9077 4320
rect 1842 3840 2158 3841
rect 1842 3776 1848 3840
rect 1912 3776 1928 3840
rect 1992 3776 2008 3840
rect 2072 3776 2088 3840
rect 2152 3776 2158 3840
rect 1842 3775 2158 3776
rect 3819 3840 4135 3841
rect 3819 3776 3825 3840
rect 3889 3776 3905 3840
rect 3969 3776 3985 3840
rect 4049 3776 4065 3840
rect 4129 3776 4135 3840
rect 3819 3775 4135 3776
rect 5796 3840 6112 3841
rect 5796 3776 5802 3840
rect 5866 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6112 3840
rect 5796 3775 6112 3776
rect 7773 3840 8089 3841
rect 7773 3776 7779 3840
rect 7843 3776 7859 3840
rect 7923 3776 7939 3840
rect 8003 3776 8019 3840
rect 8083 3776 8089 3840
rect 7773 3775 8089 3776
rect 2830 3296 3146 3297
rect 2830 3232 2836 3296
rect 2900 3232 2916 3296
rect 2980 3232 2996 3296
rect 3060 3232 3076 3296
rect 3140 3232 3146 3296
rect 2830 3231 3146 3232
rect 4807 3296 5123 3297
rect 4807 3232 4813 3296
rect 4877 3232 4893 3296
rect 4957 3232 4973 3296
rect 5037 3232 5053 3296
rect 5117 3232 5123 3296
rect 4807 3231 5123 3232
rect 6784 3296 7100 3297
rect 6784 3232 6790 3296
rect 6854 3232 6870 3296
rect 6934 3232 6950 3296
rect 7014 3232 7030 3296
rect 7094 3232 7100 3296
rect 6784 3231 7100 3232
rect 8761 3296 9077 3297
rect 8761 3232 8767 3296
rect 8831 3232 8847 3296
rect 8911 3232 8927 3296
rect 8991 3232 9007 3296
rect 9071 3232 9077 3296
rect 8761 3231 9077 3232
rect 7649 3090 7715 3093
rect 9600 3090 10000 3120
rect 7649 3088 10000 3090
rect 7649 3032 7654 3088
rect 7710 3032 10000 3088
rect 7649 3030 10000 3032
rect 7649 3027 7715 3030
rect 9600 3000 10000 3030
rect 1842 2752 2158 2753
rect 1842 2688 1848 2752
rect 1912 2688 1928 2752
rect 1992 2688 2008 2752
rect 2072 2688 2088 2752
rect 2152 2688 2158 2752
rect 1842 2687 2158 2688
rect 3819 2752 4135 2753
rect 3819 2688 3825 2752
rect 3889 2688 3905 2752
rect 3969 2688 3985 2752
rect 4049 2688 4065 2752
rect 4129 2688 4135 2752
rect 3819 2687 4135 2688
rect 5796 2752 6112 2753
rect 5796 2688 5802 2752
rect 5866 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6112 2752
rect 5796 2687 6112 2688
rect 7773 2752 8089 2753
rect 7773 2688 7779 2752
rect 7843 2688 7859 2752
rect 7923 2688 7939 2752
rect 8003 2688 8019 2752
rect 8083 2688 8089 2752
rect 7773 2687 8089 2688
rect 2830 2208 3146 2209
rect 2830 2144 2836 2208
rect 2900 2144 2916 2208
rect 2980 2144 2996 2208
rect 3060 2144 3076 2208
rect 3140 2144 3146 2208
rect 2830 2143 3146 2144
rect 4807 2208 5123 2209
rect 4807 2144 4813 2208
rect 4877 2144 4893 2208
rect 4957 2144 4973 2208
rect 5037 2144 5053 2208
rect 5117 2144 5123 2208
rect 4807 2143 5123 2144
rect 6784 2208 7100 2209
rect 6784 2144 6790 2208
rect 6854 2144 6870 2208
rect 6934 2144 6950 2208
rect 7014 2144 7030 2208
rect 7094 2144 7100 2208
rect 6784 2143 7100 2144
rect 8761 2208 9077 2209
rect 8761 2144 8767 2208
rect 8831 2144 8847 2208
rect 8911 2144 8927 2208
rect 8991 2144 9007 2208
rect 9071 2144 9077 2208
rect 8761 2143 9077 2144
rect 1842 1664 2158 1665
rect 1842 1600 1848 1664
rect 1912 1600 1928 1664
rect 1992 1600 2008 1664
rect 2072 1600 2088 1664
rect 2152 1600 2158 1664
rect 1842 1599 2158 1600
rect 3819 1664 4135 1665
rect 3819 1600 3825 1664
rect 3889 1600 3905 1664
rect 3969 1600 3985 1664
rect 4049 1600 4065 1664
rect 4129 1600 4135 1664
rect 3819 1599 4135 1600
rect 5796 1664 6112 1665
rect 5796 1600 5802 1664
rect 5866 1600 5882 1664
rect 5946 1600 5962 1664
rect 6026 1600 6042 1664
rect 6106 1600 6112 1664
rect 5796 1599 6112 1600
rect 7773 1664 8089 1665
rect 7773 1600 7779 1664
rect 7843 1600 7859 1664
rect 7923 1600 7939 1664
rect 8003 1600 8019 1664
rect 8083 1600 8089 1664
rect 7773 1599 8089 1600
rect 9305 1186 9371 1189
rect 9600 1186 10000 1216
rect 9305 1184 10000 1186
rect 9305 1128 9310 1184
rect 9366 1128 10000 1184
rect 9305 1126 10000 1128
rect 9305 1123 9371 1126
rect 2830 1120 3146 1121
rect 2830 1056 2836 1120
rect 2900 1056 2916 1120
rect 2980 1056 2996 1120
rect 3060 1056 3076 1120
rect 3140 1056 3146 1120
rect 2830 1055 3146 1056
rect 4807 1120 5123 1121
rect 4807 1056 4813 1120
rect 4877 1056 4893 1120
rect 4957 1056 4973 1120
rect 5037 1056 5053 1120
rect 5117 1056 5123 1120
rect 4807 1055 5123 1056
rect 6784 1120 7100 1121
rect 6784 1056 6790 1120
rect 6854 1056 6870 1120
rect 6934 1056 6950 1120
rect 7014 1056 7030 1120
rect 7094 1056 7100 1120
rect 6784 1055 7100 1056
rect 8761 1120 9077 1121
rect 8761 1056 8767 1120
rect 8831 1056 8847 1120
rect 8911 1056 8927 1120
rect 8991 1056 9007 1120
rect 9071 1056 9077 1120
rect 9600 1096 10000 1126
rect 8761 1055 9077 1056
<< via3 >>
rect 1848 14716 1912 14720
rect 1848 14660 1852 14716
rect 1852 14660 1908 14716
rect 1908 14660 1912 14716
rect 1848 14656 1912 14660
rect 1928 14716 1992 14720
rect 1928 14660 1932 14716
rect 1932 14660 1988 14716
rect 1988 14660 1992 14716
rect 1928 14656 1992 14660
rect 2008 14716 2072 14720
rect 2008 14660 2012 14716
rect 2012 14660 2068 14716
rect 2068 14660 2072 14716
rect 2008 14656 2072 14660
rect 2088 14716 2152 14720
rect 2088 14660 2092 14716
rect 2092 14660 2148 14716
rect 2148 14660 2152 14716
rect 2088 14656 2152 14660
rect 3825 14716 3889 14720
rect 3825 14660 3829 14716
rect 3829 14660 3885 14716
rect 3885 14660 3889 14716
rect 3825 14656 3889 14660
rect 3905 14716 3969 14720
rect 3905 14660 3909 14716
rect 3909 14660 3965 14716
rect 3965 14660 3969 14716
rect 3905 14656 3969 14660
rect 3985 14716 4049 14720
rect 3985 14660 3989 14716
rect 3989 14660 4045 14716
rect 4045 14660 4049 14716
rect 3985 14656 4049 14660
rect 4065 14716 4129 14720
rect 4065 14660 4069 14716
rect 4069 14660 4125 14716
rect 4125 14660 4129 14716
rect 4065 14656 4129 14660
rect 5802 14716 5866 14720
rect 5802 14660 5806 14716
rect 5806 14660 5862 14716
rect 5862 14660 5866 14716
rect 5802 14656 5866 14660
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 7779 14716 7843 14720
rect 7779 14660 7783 14716
rect 7783 14660 7839 14716
rect 7839 14660 7843 14716
rect 7779 14656 7843 14660
rect 7859 14716 7923 14720
rect 7859 14660 7863 14716
rect 7863 14660 7919 14716
rect 7919 14660 7923 14716
rect 7859 14656 7923 14660
rect 7939 14716 8003 14720
rect 7939 14660 7943 14716
rect 7943 14660 7999 14716
rect 7999 14660 8003 14716
rect 7939 14656 8003 14660
rect 8019 14716 8083 14720
rect 8019 14660 8023 14716
rect 8023 14660 8079 14716
rect 8079 14660 8083 14716
rect 8019 14656 8083 14660
rect 2836 14172 2900 14176
rect 2836 14116 2840 14172
rect 2840 14116 2896 14172
rect 2896 14116 2900 14172
rect 2836 14112 2900 14116
rect 2916 14172 2980 14176
rect 2916 14116 2920 14172
rect 2920 14116 2976 14172
rect 2976 14116 2980 14172
rect 2916 14112 2980 14116
rect 2996 14172 3060 14176
rect 2996 14116 3000 14172
rect 3000 14116 3056 14172
rect 3056 14116 3060 14172
rect 2996 14112 3060 14116
rect 3076 14172 3140 14176
rect 3076 14116 3080 14172
rect 3080 14116 3136 14172
rect 3136 14116 3140 14172
rect 3076 14112 3140 14116
rect 4813 14172 4877 14176
rect 4813 14116 4817 14172
rect 4817 14116 4873 14172
rect 4873 14116 4877 14172
rect 4813 14112 4877 14116
rect 4893 14172 4957 14176
rect 4893 14116 4897 14172
rect 4897 14116 4953 14172
rect 4953 14116 4957 14172
rect 4893 14112 4957 14116
rect 4973 14172 5037 14176
rect 4973 14116 4977 14172
rect 4977 14116 5033 14172
rect 5033 14116 5037 14172
rect 4973 14112 5037 14116
rect 5053 14172 5117 14176
rect 5053 14116 5057 14172
rect 5057 14116 5113 14172
rect 5113 14116 5117 14172
rect 5053 14112 5117 14116
rect 6790 14172 6854 14176
rect 6790 14116 6794 14172
rect 6794 14116 6850 14172
rect 6850 14116 6854 14172
rect 6790 14112 6854 14116
rect 6870 14172 6934 14176
rect 6870 14116 6874 14172
rect 6874 14116 6930 14172
rect 6930 14116 6934 14172
rect 6870 14112 6934 14116
rect 6950 14172 7014 14176
rect 6950 14116 6954 14172
rect 6954 14116 7010 14172
rect 7010 14116 7014 14172
rect 6950 14112 7014 14116
rect 7030 14172 7094 14176
rect 7030 14116 7034 14172
rect 7034 14116 7090 14172
rect 7090 14116 7094 14172
rect 7030 14112 7094 14116
rect 8767 14172 8831 14176
rect 8767 14116 8771 14172
rect 8771 14116 8827 14172
rect 8827 14116 8831 14172
rect 8767 14112 8831 14116
rect 8847 14172 8911 14176
rect 8847 14116 8851 14172
rect 8851 14116 8907 14172
rect 8907 14116 8911 14172
rect 8847 14112 8911 14116
rect 8927 14172 8991 14176
rect 8927 14116 8931 14172
rect 8931 14116 8987 14172
rect 8987 14116 8991 14172
rect 8927 14112 8991 14116
rect 9007 14172 9071 14176
rect 9007 14116 9011 14172
rect 9011 14116 9067 14172
rect 9067 14116 9071 14172
rect 9007 14112 9071 14116
rect 1848 13628 1912 13632
rect 1848 13572 1852 13628
rect 1852 13572 1908 13628
rect 1908 13572 1912 13628
rect 1848 13568 1912 13572
rect 1928 13628 1992 13632
rect 1928 13572 1932 13628
rect 1932 13572 1988 13628
rect 1988 13572 1992 13628
rect 1928 13568 1992 13572
rect 2008 13628 2072 13632
rect 2008 13572 2012 13628
rect 2012 13572 2068 13628
rect 2068 13572 2072 13628
rect 2008 13568 2072 13572
rect 2088 13628 2152 13632
rect 2088 13572 2092 13628
rect 2092 13572 2148 13628
rect 2148 13572 2152 13628
rect 2088 13568 2152 13572
rect 3825 13628 3889 13632
rect 3825 13572 3829 13628
rect 3829 13572 3885 13628
rect 3885 13572 3889 13628
rect 3825 13568 3889 13572
rect 3905 13628 3969 13632
rect 3905 13572 3909 13628
rect 3909 13572 3965 13628
rect 3965 13572 3969 13628
rect 3905 13568 3969 13572
rect 3985 13628 4049 13632
rect 3985 13572 3989 13628
rect 3989 13572 4045 13628
rect 4045 13572 4049 13628
rect 3985 13568 4049 13572
rect 4065 13628 4129 13632
rect 4065 13572 4069 13628
rect 4069 13572 4125 13628
rect 4125 13572 4129 13628
rect 4065 13568 4129 13572
rect 5802 13628 5866 13632
rect 5802 13572 5806 13628
rect 5806 13572 5862 13628
rect 5862 13572 5866 13628
rect 5802 13568 5866 13572
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 7779 13628 7843 13632
rect 7779 13572 7783 13628
rect 7783 13572 7839 13628
rect 7839 13572 7843 13628
rect 7779 13568 7843 13572
rect 7859 13628 7923 13632
rect 7859 13572 7863 13628
rect 7863 13572 7919 13628
rect 7919 13572 7923 13628
rect 7859 13568 7923 13572
rect 7939 13628 8003 13632
rect 7939 13572 7943 13628
rect 7943 13572 7999 13628
rect 7999 13572 8003 13628
rect 7939 13568 8003 13572
rect 8019 13628 8083 13632
rect 8019 13572 8023 13628
rect 8023 13572 8079 13628
rect 8079 13572 8083 13628
rect 8019 13568 8083 13572
rect 2836 13084 2900 13088
rect 2836 13028 2840 13084
rect 2840 13028 2896 13084
rect 2896 13028 2900 13084
rect 2836 13024 2900 13028
rect 2916 13084 2980 13088
rect 2916 13028 2920 13084
rect 2920 13028 2976 13084
rect 2976 13028 2980 13084
rect 2916 13024 2980 13028
rect 2996 13084 3060 13088
rect 2996 13028 3000 13084
rect 3000 13028 3056 13084
rect 3056 13028 3060 13084
rect 2996 13024 3060 13028
rect 3076 13084 3140 13088
rect 3076 13028 3080 13084
rect 3080 13028 3136 13084
rect 3136 13028 3140 13084
rect 3076 13024 3140 13028
rect 4813 13084 4877 13088
rect 4813 13028 4817 13084
rect 4817 13028 4873 13084
rect 4873 13028 4877 13084
rect 4813 13024 4877 13028
rect 4893 13084 4957 13088
rect 4893 13028 4897 13084
rect 4897 13028 4953 13084
rect 4953 13028 4957 13084
rect 4893 13024 4957 13028
rect 4973 13084 5037 13088
rect 4973 13028 4977 13084
rect 4977 13028 5033 13084
rect 5033 13028 5037 13084
rect 4973 13024 5037 13028
rect 5053 13084 5117 13088
rect 5053 13028 5057 13084
rect 5057 13028 5113 13084
rect 5113 13028 5117 13084
rect 5053 13024 5117 13028
rect 6790 13084 6854 13088
rect 6790 13028 6794 13084
rect 6794 13028 6850 13084
rect 6850 13028 6854 13084
rect 6790 13024 6854 13028
rect 6870 13084 6934 13088
rect 6870 13028 6874 13084
rect 6874 13028 6930 13084
rect 6930 13028 6934 13084
rect 6870 13024 6934 13028
rect 6950 13084 7014 13088
rect 6950 13028 6954 13084
rect 6954 13028 7010 13084
rect 7010 13028 7014 13084
rect 6950 13024 7014 13028
rect 7030 13084 7094 13088
rect 7030 13028 7034 13084
rect 7034 13028 7090 13084
rect 7090 13028 7094 13084
rect 7030 13024 7094 13028
rect 8767 13084 8831 13088
rect 8767 13028 8771 13084
rect 8771 13028 8827 13084
rect 8827 13028 8831 13084
rect 8767 13024 8831 13028
rect 8847 13084 8911 13088
rect 8847 13028 8851 13084
rect 8851 13028 8907 13084
rect 8907 13028 8911 13084
rect 8847 13024 8911 13028
rect 8927 13084 8991 13088
rect 8927 13028 8931 13084
rect 8931 13028 8987 13084
rect 8987 13028 8991 13084
rect 8927 13024 8991 13028
rect 9007 13084 9071 13088
rect 9007 13028 9011 13084
rect 9011 13028 9067 13084
rect 9067 13028 9071 13084
rect 9007 13024 9071 13028
rect 1848 12540 1912 12544
rect 1848 12484 1852 12540
rect 1852 12484 1908 12540
rect 1908 12484 1912 12540
rect 1848 12480 1912 12484
rect 1928 12540 1992 12544
rect 1928 12484 1932 12540
rect 1932 12484 1988 12540
rect 1988 12484 1992 12540
rect 1928 12480 1992 12484
rect 2008 12540 2072 12544
rect 2008 12484 2012 12540
rect 2012 12484 2068 12540
rect 2068 12484 2072 12540
rect 2008 12480 2072 12484
rect 2088 12540 2152 12544
rect 2088 12484 2092 12540
rect 2092 12484 2148 12540
rect 2148 12484 2152 12540
rect 2088 12480 2152 12484
rect 3825 12540 3889 12544
rect 3825 12484 3829 12540
rect 3829 12484 3885 12540
rect 3885 12484 3889 12540
rect 3825 12480 3889 12484
rect 3905 12540 3969 12544
rect 3905 12484 3909 12540
rect 3909 12484 3965 12540
rect 3965 12484 3969 12540
rect 3905 12480 3969 12484
rect 3985 12540 4049 12544
rect 3985 12484 3989 12540
rect 3989 12484 4045 12540
rect 4045 12484 4049 12540
rect 3985 12480 4049 12484
rect 4065 12540 4129 12544
rect 4065 12484 4069 12540
rect 4069 12484 4125 12540
rect 4125 12484 4129 12540
rect 4065 12480 4129 12484
rect 5802 12540 5866 12544
rect 5802 12484 5806 12540
rect 5806 12484 5862 12540
rect 5862 12484 5866 12540
rect 5802 12480 5866 12484
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 7779 12540 7843 12544
rect 7779 12484 7783 12540
rect 7783 12484 7839 12540
rect 7839 12484 7843 12540
rect 7779 12480 7843 12484
rect 7859 12540 7923 12544
rect 7859 12484 7863 12540
rect 7863 12484 7919 12540
rect 7919 12484 7923 12540
rect 7859 12480 7923 12484
rect 7939 12540 8003 12544
rect 7939 12484 7943 12540
rect 7943 12484 7999 12540
rect 7999 12484 8003 12540
rect 7939 12480 8003 12484
rect 8019 12540 8083 12544
rect 8019 12484 8023 12540
rect 8023 12484 8079 12540
rect 8079 12484 8083 12540
rect 8019 12480 8083 12484
rect 2836 11996 2900 12000
rect 2836 11940 2840 11996
rect 2840 11940 2896 11996
rect 2896 11940 2900 11996
rect 2836 11936 2900 11940
rect 2916 11996 2980 12000
rect 2916 11940 2920 11996
rect 2920 11940 2976 11996
rect 2976 11940 2980 11996
rect 2916 11936 2980 11940
rect 2996 11996 3060 12000
rect 2996 11940 3000 11996
rect 3000 11940 3056 11996
rect 3056 11940 3060 11996
rect 2996 11936 3060 11940
rect 3076 11996 3140 12000
rect 3076 11940 3080 11996
rect 3080 11940 3136 11996
rect 3136 11940 3140 11996
rect 3076 11936 3140 11940
rect 4813 11996 4877 12000
rect 4813 11940 4817 11996
rect 4817 11940 4873 11996
rect 4873 11940 4877 11996
rect 4813 11936 4877 11940
rect 4893 11996 4957 12000
rect 4893 11940 4897 11996
rect 4897 11940 4953 11996
rect 4953 11940 4957 11996
rect 4893 11936 4957 11940
rect 4973 11996 5037 12000
rect 4973 11940 4977 11996
rect 4977 11940 5033 11996
rect 5033 11940 5037 11996
rect 4973 11936 5037 11940
rect 5053 11996 5117 12000
rect 5053 11940 5057 11996
rect 5057 11940 5113 11996
rect 5113 11940 5117 11996
rect 5053 11936 5117 11940
rect 6790 11996 6854 12000
rect 6790 11940 6794 11996
rect 6794 11940 6850 11996
rect 6850 11940 6854 11996
rect 6790 11936 6854 11940
rect 6870 11996 6934 12000
rect 6870 11940 6874 11996
rect 6874 11940 6930 11996
rect 6930 11940 6934 11996
rect 6870 11936 6934 11940
rect 6950 11996 7014 12000
rect 6950 11940 6954 11996
rect 6954 11940 7010 11996
rect 7010 11940 7014 11996
rect 6950 11936 7014 11940
rect 7030 11996 7094 12000
rect 7030 11940 7034 11996
rect 7034 11940 7090 11996
rect 7090 11940 7094 11996
rect 7030 11936 7094 11940
rect 8767 11996 8831 12000
rect 8767 11940 8771 11996
rect 8771 11940 8827 11996
rect 8827 11940 8831 11996
rect 8767 11936 8831 11940
rect 8847 11996 8911 12000
rect 8847 11940 8851 11996
rect 8851 11940 8907 11996
rect 8907 11940 8911 11996
rect 8847 11936 8911 11940
rect 8927 11996 8991 12000
rect 8927 11940 8931 11996
rect 8931 11940 8987 11996
rect 8987 11940 8991 11996
rect 8927 11936 8991 11940
rect 9007 11996 9071 12000
rect 9007 11940 9011 11996
rect 9011 11940 9067 11996
rect 9067 11940 9071 11996
rect 9007 11936 9071 11940
rect 1848 11452 1912 11456
rect 1848 11396 1852 11452
rect 1852 11396 1908 11452
rect 1908 11396 1912 11452
rect 1848 11392 1912 11396
rect 1928 11452 1992 11456
rect 1928 11396 1932 11452
rect 1932 11396 1988 11452
rect 1988 11396 1992 11452
rect 1928 11392 1992 11396
rect 2008 11452 2072 11456
rect 2008 11396 2012 11452
rect 2012 11396 2068 11452
rect 2068 11396 2072 11452
rect 2008 11392 2072 11396
rect 2088 11452 2152 11456
rect 2088 11396 2092 11452
rect 2092 11396 2148 11452
rect 2148 11396 2152 11452
rect 2088 11392 2152 11396
rect 3825 11452 3889 11456
rect 3825 11396 3829 11452
rect 3829 11396 3885 11452
rect 3885 11396 3889 11452
rect 3825 11392 3889 11396
rect 3905 11452 3969 11456
rect 3905 11396 3909 11452
rect 3909 11396 3965 11452
rect 3965 11396 3969 11452
rect 3905 11392 3969 11396
rect 3985 11452 4049 11456
rect 3985 11396 3989 11452
rect 3989 11396 4045 11452
rect 4045 11396 4049 11452
rect 3985 11392 4049 11396
rect 4065 11452 4129 11456
rect 4065 11396 4069 11452
rect 4069 11396 4125 11452
rect 4125 11396 4129 11452
rect 4065 11392 4129 11396
rect 5802 11452 5866 11456
rect 5802 11396 5806 11452
rect 5806 11396 5862 11452
rect 5862 11396 5866 11452
rect 5802 11392 5866 11396
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 7779 11452 7843 11456
rect 7779 11396 7783 11452
rect 7783 11396 7839 11452
rect 7839 11396 7843 11452
rect 7779 11392 7843 11396
rect 7859 11452 7923 11456
rect 7859 11396 7863 11452
rect 7863 11396 7919 11452
rect 7919 11396 7923 11452
rect 7859 11392 7923 11396
rect 7939 11452 8003 11456
rect 7939 11396 7943 11452
rect 7943 11396 7999 11452
rect 7999 11396 8003 11452
rect 7939 11392 8003 11396
rect 8019 11452 8083 11456
rect 8019 11396 8023 11452
rect 8023 11396 8079 11452
rect 8079 11396 8083 11452
rect 8019 11392 8083 11396
rect 2836 10908 2900 10912
rect 2836 10852 2840 10908
rect 2840 10852 2896 10908
rect 2896 10852 2900 10908
rect 2836 10848 2900 10852
rect 2916 10908 2980 10912
rect 2916 10852 2920 10908
rect 2920 10852 2976 10908
rect 2976 10852 2980 10908
rect 2916 10848 2980 10852
rect 2996 10908 3060 10912
rect 2996 10852 3000 10908
rect 3000 10852 3056 10908
rect 3056 10852 3060 10908
rect 2996 10848 3060 10852
rect 3076 10908 3140 10912
rect 3076 10852 3080 10908
rect 3080 10852 3136 10908
rect 3136 10852 3140 10908
rect 3076 10848 3140 10852
rect 4813 10908 4877 10912
rect 4813 10852 4817 10908
rect 4817 10852 4873 10908
rect 4873 10852 4877 10908
rect 4813 10848 4877 10852
rect 4893 10908 4957 10912
rect 4893 10852 4897 10908
rect 4897 10852 4953 10908
rect 4953 10852 4957 10908
rect 4893 10848 4957 10852
rect 4973 10908 5037 10912
rect 4973 10852 4977 10908
rect 4977 10852 5033 10908
rect 5033 10852 5037 10908
rect 4973 10848 5037 10852
rect 5053 10908 5117 10912
rect 5053 10852 5057 10908
rect 5057 10852 5113 10908
rect 5113 10852 5117 10908
rect 5053 10848 5117 10852
rect 6790 10908 6854 10912
rect 6790 10852 6794 10908
rect 6794 10852 6850 10908
rect 6850 10852 6854 10908
rect 6790 10848 6854 10852
rect 6870 10908 6934 10912
rect 6870 10852 6874 10908
rect 6874 10852 6930 10908
rect 6930 10852 6934 10908
rect 6870 10848 6934 10852
rect 6950 10908 7014 10912
rect 6950 10852 6954 10908
rect 6954 10852 7010 10908
rect 7010 10852 7014 10908
rect 6950 10848 7014 10852
rect 7030 10908 7094 10912
rect 7030 10852 7034 10908
rect 7034 10852 7090 10908
rect 7090 10852 7094 10908
rect 7030 10848 7094 10852
rect 8767 10908 8831 10912
rect 8767 10852 8771 10908
rect 8771 10852 8827 10908
rect 8827 10852 8831 10908
rect 8767 10848 8831 10852
rect 8847 10908 8911 10912
rect 8847 10852 8851 10908
rect 8851 10852 8907 10908
rect 8907 10852 8911 10908
rect 8847 10848 8911 10852
rect 8927 10908 8991 10912
rect 8927 10852 8931 10908
rect 8931 10852 8987 10908
rect 8987 10852 8991 10908
rect 8927 10848 8991 10852
rect 9007 10908 9071 10912
rect 9007 10852 9011 10908
rect 9011 10852 9067 10908
rect 9067 10852 9071 10908
rect 9007 10848 9071 10852
rect 1848 10364 1912 10368
rect 1848 10308 1852 10364
rect 1852 10308 1908 10364
rect 1908 10308 1912 10364
rect 1848 10304 1912 10308
rect 1928 10364 1992 10368
rect 1928 10308 1932 10364
rect 1932 10308 1988 10364
rect 1988 10308 1992 10364
rect 1928 10304 1992 10308
rect 2008 10364 2072 10368
rect 2008 10308 2012 10364
rect 2012 10308 2068 10364
rect 2068 10308 2072 10364
rect 2008 10304 2072 10308
rect 2088 10364 2152 10368
rect 2088 10308 2092 10364
rect 2092 10308 2148 10364
rect 2148 10308 2152 10364
rect 2088 10304 2152 10308
rect 3825 10364 3889 10368
rect 3825 10308 3829 10364
rect 3829 10308 3885 10364
rect 3885 10308 3889 10364
rect 3825 10304 3889 10308
rect 3905 10364 3969 10368
rect 3905 10308 3909 10364
rect 3909 10308 3965 10364
rect 3965 10308 3969 10364
rect 3905 10304 3969 10308
rect 3985 10364 4049 10368
rect 3985 10308 3989 10364
rect 3989 10308 4045 10364
rect 4045 10308 4049 10364
rect 3985 10304 4049 10308
rect 4065 10364 4129 10368
rect 4065 10308 4069 10364
rect 4069 10308 4125 10364
rect 4125 10308 4129 10364
rect 4065 10304 4129 10308
rect 5802 10364 5866 10368
rect 5802 10308 5806 10364
rect 5806 10308 5862 10364
rect 5862 10308 5866 10364
rect 5802 10304 5866 10308
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 7779 10364 7843 10368
rect 7779 10308 7783 10364
rect 7783 10308 7839 10364
rect 7839 10308 7843 10364
rect 7779 10304 7843 10308
rect 7859 10364 7923 10368
rect 7859 10308 7863 10364
rect 7863 10308 7919 10364
rect 7919 10308 7923 10364
rect 7859 10304 7923 10308
rect 7939 10364 8003 10368
rect 7939 10308 7943 10364
rect 7943 10308 7999 10364
rect 7999 10308 8003 10364
rect 7939 10304 8003 10308
rect 8019 10364 8083 10368
rect 8019 10308 8023 10364
rect 8023 10308 8079 10364
rect 8079 10308 8083 10364
rect 8019 10304 8083 10308
rect 2836 9820 2900 9824
rect 2836 9764 2840 9820
rect 2840 9764 2896 9820
rect 2896 9764 2900 9820
rect 2836 9760 2900 9764
rect 2916 9820 2980 9824
rect 2916 9764 2920 9820
rect 2920 9764 2976 9820
rect 2976 9764 2980 9820
rect 2916 9760 2980 9764
rect 2996 9820 3060 9824
rect 2996 9764 3000 9820
rect 3000 9764 3056 9820
rect 3056 9764 3060 9820
rect 2996 9760 3060 9764
rect 3076 9820 3140 9824
rect 3076 9764 3080 9820
rect 3080 9764 3136 9820
rect 3136 9764 3140 9820
rect 3076 9760 3140 9764
rect 4813 9820 4877 9824
rect 4813 9764 4817 9820
rect 4817 9764 4873 9820
rect 4873 9764 4877 9820
rect 4813 9760 4877 9764
rect 4893 9820 4957 9824
rect 4893 9764 4897 9820
rect 4897 9764 4953 9820
rect 4953 9764 4957 9820
rect 4893 9760 4957 9764
rect 4973 9820 5037 9824
rect 4973 9764 4977 9820
rect 4977 9764 5033 9820
rect 5033 9764 5037 9820
rect 4973 9760 5037 9764
rect 5053 9820 5117 9824
rect 5053 9764 5057 9820
rect 5057 9764 5113 9820
rect 5113 9764 5117 9820
rect 5053 9760 5117 9764
rect 6790 9820 6854 9824
rect 6790 9764 6794 9820
rect 6794 9764 6850 9820
rect 6850 9764 6854 9820
rect 6790 9760 6854 9764
rect 6870 9820 6934 9824
rect 6870 9764 6874 9820
rect 6874 9764 6930 9820
rect 6930 9764 6934 9820
rect 6870 9760 6934 9764
rect 6950 9820 7014 9824
rect 6950 9764 6954 9820
rect 6954 9764 7010 9820
rect 7010 9764 7014 9820
rect 6950 9760 7014 9764
rect 7030 9820 7094 9824
rect 7030 9764 7034 9820
rect 7034 9764 7090 9820
rect 7090 9764 7094 9820
rect 7030 9760 7094 9764
rect 8767 9820 8831 9824
rect 8767 9764 8771 9820
rect 8771 9764 8827 9820
rect 8827 9764 8831 9820
rect 8767 9760 8831 9764
rect 8847 9820 8911 9824
rect 8847 9764 8851 9820
rect 8851 9764 8907 9820
rect 8907 9764 8911 9820
rect 8847 9760 8911 9764
rect 8927 9820 8991 9824
rect 8927 9764 8931 9820
rect 8931 9764 8987 9820
rect 8987 9764 8991 9820
rect 8927 9760 8991 9764
rect 9007 9820 9071 9824
rect 9007 9764 9011 9820
rect 9011 9764 9067 9820
rect 9067 9764 9071 9820
rect 9007 9760 9071 9764
rect 1848 9276 1912 9280
rect 1848 9220 1852 9276
rect 1852 9220 1908 9276
rect 1908 9220 1912 9276
rect 1848 9216 1912 9220
rect 1928 9276 1992 9280
rect 1928 9220 1932 9276
rect 1932 9220 1988 9276
rect 1988 9220 1992 9276
rect 1928 9216 1992 9220
rect 2008 9276 2072 9280
rect 2008 9220 2012 9276
rect 2012 9220 2068 9276
rect 2068 9220 2072 9276
rect 2008 9216 2072 9220
rect 2088 9276 2152 9280
rect 2088 9220 2092 9276
rect 2092 9220 2148 9276
rect 2148 9220 2152 9276
rect 2088 9216 2152 9220
rect 3825 9276 3889 9280
rect 3825 9220 3829 9276
rect 3829 9220 3885 9276
rect 3885 9220 3889 9276
rect 3825 9216 3889 9220
rect 3905 9276 3969 9280
rect 3905 9220 3909 9276
rect 3909 9220 3965 9276
rect 3965 9220 3969 9276
rect 3905 9216 3969 9220
rect 3985 9276 4049 9280
rect 3985 9220 3989 9276
rect 3989 9220 4045 9276
rect 4045 9220 4049 9276
rect 3985 9216 4049 9220
rect 4065 9276 4129 9280
rect 4065 9220 4069 9276
rect 4069 9220 4125 9276
rect 4125 9220 4129 9276
rect 4065 9216 4129 9220
rect 5802 9276 5866 9280
rect 5802 9220 5806 9276
rect 5806 9220 5862 9276
rect 5862 9220 5866 9276
rect 5802 9216 5866 9220
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 7779 9276 7843 9280
rect 7779 9220 7783 9276
rect 7783 9220 7839 9276
rect 7839 9220 7843 9276
rect 7779 9216 7843 9220
rect 7859 9276 7923 9280
rect 7859 9220 7863 9276
rect 7863 9220 7919 9276
rect 7919 9220 7923 9276
rect 7859 9216 7923 9220
rect 7939 9276 8003 9280
rect 7939 9220 7943 9276
rect 7943 9220 7999 9276
rect 7999 9220 8003 9276
rect 7939 9216 8003 9220
rect 8019 9276 8083 9280
rect 8019 9220 8023 9276
rect 8023 9220 8079 9276
rect 8079 9220 8083 9276
rect 8019 9216 8083 9220
rect 2836 8732 2900 8736
rect 2836 8676 2840 8732
rect 2840 8676 2896 8732
rect 2896 8676 2900 8732
rect 2836 8672 2900 8676
rect 2916 8732 2980 8736
rect 2916 8676 2920 8732
rect 2920 8676 2976 8732
rect 2976 8676 2980 8732
rect 2916 8672 2980 8676
rect 2996 8732 3060 8736
rect 2996 8676 3000 8732
rect 3000 8676 3056 8732
rect 3056 8676 3060 8732
rect 2996 8672 3060 8676
rect 3076 8732 3140 8736
rect 3076 8676 3080 8732
rect 3080 8676 3136 8732
rect 3136 8676 3140 8732
rect 3076 8672 3140 8676
rect 4813 8732 4877 8736
rect 4813 8676 4817 8732
rect 4817 8676 4873 8732
rect 4873 8676 4877 8732
rect 4813 8672 4877 8676
rect 4893 8732 4957 8736
rect 4893 8676 4897 8732
rect 4897 8676 4953 8732
rect 4953 8676 4957 8732
rect 4893 8672 4957 8676
rect 4973 8732 5037 8736
rect 4973 8676 4977 8732
rect 4977 8676 5033 8732
rect 5033 8676 5037 8732
rect 4973 8672 5037 8676
rect 5053 8732 5117 8736
rect 5053 8676 5057 8732
rect 5057 8676 5113 8732
rect 5113 8676 5117 8732
rect 5053 8672 5117 8676
rect 6790 8732 6854 8736
rect 6790 8676 6794 8732
rect 6794 8676 6850 8732
rect 6850 8676 6854 8732
rect 6790 8672 6854 8676
rect 6870 8732 6934 8736
rect 6870 8676 6874 8732
rect 6874 8676 6930 8732
rect 6930 8676 6934 8732
rect 6870 8672 6934 8676
rect 6950 8732 7014 8736
rect 6950 8676 6954 8732
rect 6954 8676 7010 8732
rect 7010 8676 7014 8732
rect 6950 8672 7014 8676
rect 7030 8732 7094 8736
rect 7030 8676 7034 8732
rect 7034 8676 7090 8732
rect 7090 8676 7094 8732
rect 7030 8672 7094 8676
rect 8767 8732 8831 8736
rect 8767 8676 8771 8732
rect 8771 8676 8827 8732
rect 8827 8676 8831 8732
rect 8767 8672 8831 8676
rect 8847 8732 8911 8736
rect 8847 8676 8851 8732
rect 8851 8676 8907 8732
rect 8907 8676 8911 8732
rect 8847 8672 8911 8676
rect 8927 8732 8991 8736
rect 8927 8676 8931 8732
rect 8931 8676 8987 8732
rect 8987 8676 8991 8732
rect 8927 8672 8991 8676
rect 9007 8732 9071 8736
rect 9007 8676 9011 8732
rect 9011 8676 9067 8732
rect 9067 8676 9071 8732
rect 9007 8672 9071 8676
rect 1848 8188 1912 8192
rect 1848 8132 1852 8188
rect 1852 8132 1908 8188
rect 1908 8132 1912 8188
rect 1848 8128 1912 8132
rect 1928 8188 1992 8192
rect 1928 8132 1932 8188
rect 1932 8132 1988 8188
rect 1988 8132 1992 8188
rect 1928 8128 1992 8132
rect 2008 8188 2072 8192
rect 2008 8132 2012 8188
rect 2012 8132 2068 8188
rect 2068 8132 2072 8188
rect 2008 8128 2072 8132
rect 2088 8188 2152 8192
rect 2088 8132 2092 8188
rect 2092 8132 2148 8188
rect 2148 8132 2152 8188
rect 2088 8128 2152 8132
rect 3825 8188 3889 8192
rect 3825 8132 3829 8188
rect 3829 8132 3885 8188
rect 3885 8132 3889 8188
rect 3825 8128 3889 8132
rect 3905 8188 3969 8192
rect 3905 8132 3909 8188
rect 3909 8132 3965 8188
rect 3965 8132 3969 8188
rect 3905 8128 3969 8132
rect 3985 8188 4049 8192
rect 3985 8132 3989 8188
rect 3989 8132 4045 8188
rect 4045 8132 4049 8188
rect 3985 8128 4049 8132
rect 4065 8188 4129 8192
rect 4065 8132 4069 8188
rect 4069 8132 4125 8188
rect 4125 8132 4129 8188
rect 4065 8128 4129 8132
rect 5802 8188 5866 8192
rect 5802 8132 5806 8188
rect 5806 8132 5862 8188
rect 5862 8132 5866 8188
rect 5802 8128 5866 8132
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 7779 8188 7843 8192
rect 7779 8132 7783 8188
rect 7783 8132 7839 8188
rect 7839 8132 7843 8188
rect 7779 8128 7843 8132
rect 7859 8188 7923 8192
rect 7859 8132 7863 8188
rect 7863 8132 7919 8188
rect 7919 8132 7923 8188
rect 7859 8128 7923 8132
rect 7939 8188 8003 8192
rect 7939 8132 7943 8188
rect 7943 8132 7999 8188
rect 7999 8132 8003 8188
rect 7939 8128 8003 8132
rect 8019 8188 8083 8192
rect 8019 8132 8023 8188
rect 8023 8132 8079 8188
rect 8079 8132 8083 8188
rect 8019 8128 8083 8132
rect 2836 7644 2900 7648
rect 2836 7588 2840 7644
rect 2840 7588 2896 7644
rect 2896 7588 2900 7644
rect 2836 7584 2900 7588
rect 2916 7644 2980 7648
rect 2916 7588 2920 7644
rect 2920 7588 2976 7644
rect 2976 7588 2980 7644
rect 2916 7584 2980 7588
rect 2996 7644 3060 7648
rect 2996 7588 3000 7644
rect 3000 7588 3056 7644
rect 3056 7588 3060 7644
rect 2996 7584 3060 7588
rect 3076 7644 3140 7648
rect 3076 7588 3080 7644
rect 3080 7588 3136 7644
rect 3136 7588 3140 7644
rect 3076 7584 3140 7588
rect 4813 7644 4877 7648
rect 4813 7588 4817 7644
rect 4817 7588 4873 7644
rect 4873 7588 4877 7644
rect 4813 7584 4877 7588
rect 4893 7644 4957 7648
rect 4893 7588 4897 7644
rect 4897 7588 4953 7644
rect 4953 7588 4957 7644
rect 4893 7584 4957 7588
rect 4973 7644 5037 7648
rect 4973 7588 4977 7644
rect 4977 7588 5033 7644
rect 5033 7588 5037 7644
rect 4973 7584 5037 7588
rect 5053 7644 5117 7648
rect 5053 7588 5057 7644
rect 5057 7588 5113 7644
rect 5113 7588 5117 7644
rect 5053 7584 5117 7588
rect 6790 7644 6854 7648
rect 6790 7588 6794 7644
rect 6794 7588 6850 7644
rect 6850 7588 6854 7644
rect 6790 7584 6854 7588
rect 6870 7644 6934 7648
rect 6870 7588 6874 7644
rect 6874 7588 6930 7644
rect 6930 7588 6934 7644
rect 6870 7584 6934 7588
rect 6950 7644 7014 7648
rect 6950 7588 6954 7644
rect 6954 7588 7010 7644
rect 7010 7588 7014 7644
rect 6950 7584 7014 7588
rect 7030 7644 7094 7648
rect 7030 7588 7034 7644
rect 7034 7588 7090 7644
rect 7090 7588 7094 7644
rect 7030 7584 7094 7588
rect 8767 7644 8831 7648
rect 8767 7588 8771 7644
rect 8771 7588 8827 7644
rect 8827 7588 8831 7644
rect 8767 7584 8831 7588
rect 8847 7644 8911 7648
rect 8847 7588 8851 7644
rect 8851 7588 8907 7644
rect 8907 7588 8911 7644
rect 8847 7584 8911 7588
rect 8927 7644 8991 7648
rect 8927 7588 8931 7644
rect 8931 7588 8987 7644
rect 8987 7588 8991 7644
rect 8927 7584 8991 7588
rect 9007 7644 9071 7648
rect 9007 7588 9011 7644
rect 9011 7588 9067 7644
rect 9067 7588 9071 7644
rect 9007 7584 9071 7588
rect 1848 7100 1912 7104
rect 1848 7044 1852 7100
rect 1852 7044 1908 7100
rect 1908 7044 1912 7100
rect 1848 7040 1912 7044
rect 1928 7100 1992 7104
rect 1928 7044 1932 7100
rect 1932 7044 1988 7100
rect 1988 7044 1992 7100
rect 1928 7040 1992 7044
rect 2008 7100 2072 7104
rect 2008 7044 2012 7100
rect 2012 7044 2068 7100
rect 2068 7044 2072 7100
rect 2008 7040 2072 7044
rect 2088 7100 2152 7104
rect 2088 7044 2092 7100
rect 2092 7044 2148 7100
rect 2148 7044 2152 7100
rect 2088 7040 2152 7044
rect 3825 7100 3889 7104
rect 3825 7044 3829 7100
rect 3829 7044 3885 7100
rect 3885 7044 3889 7100
rect 3825 7040 3889 7044
rect 3905 7100 3969 7104
rect 3905 7044 3909 7100
rect 3909 7044 3965 7100
rect 3965 7044 3969 7100
rect 3905 7040 3969 7044
rect 3985 7100 4049 7104
rect 3985 7044 3989 7100
rect 3989 7044 4045 7100
rect 4045 7044 4049 7100
rect 3985 7040 4049 7044
rect 4065 7100 4129 7104
rect 4065 7044 4069 7100
rect 4069 7044 4125 7100
rect 4125 7044 4129 7100
rect 4065 7040 4129 7044
rect 5802 7100 5866 7104
rect 5802 7044 5806 7100
rect 5806 7044 5862 7100
rect 5862 7044 5866 7100
rect 5802 7040 5866 7044
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 7779 7100 7843 7104
rect 7779 7044 7783 7100
rect 7783 7044 7839 7100
rect 7839 7044 7843 7100
rect 7779 7040 7843 7044
rect 7859 7100 7923 7104
rect 7859 7044 7863 7100
rect 7863 7044 7919 7100
rect 7919 7044 7923 7100
rect 7859 7040 7923 7044
rect 7939 7100 8003 7104
rect 7939 7044 7943 7100
rect 7943 7044 7999 7100
rect 7999 7044 8003 7100
rect 7939 7040 8003 7044
rect 8019 7100 8083 7104
rect 8019 7044 8023 7100
rect 8023 7044 8079 7100
rect 8079 7044 8083 7100
rect 8019 7040 8083 7044
rect 2836 6556 2900 6560
rect 2836 6500 2840 6556
rect 2840 6500 2896 6556
rect 2896 6500 2900 6556
rect 2836 6496 2900 6500
rect 2916 6556 2980 6560
rect 2916 6500 2920 6556
rect 2920 6500 2976 6556
rect 2976 6500 2980 6556
rect 2916 6496 2980 6500
rect 2996 6556 3060 6560
rect 2996 6500 3000 6556
rect 3000 6500 3056 6556
rect 3056 6500 3060 6556
rect 2996 6496 3060 6500
rect 3076 6556 3140 6560
rect 3076 6500 3080 6556
rect 3080 6500 3136 6556
rect 3136 6500 3140 6556
rect 3076 6496 3140 6500
rect 4813 6556 4877 6560
rect 4813 6500 4817 6556
rect 4817 6500 4873 6556
rect 4873 6500 4877 6556
rect 4813 6496 4877 6500
rect 4893 6556 4957 6560
rect 4893 6500 4897 6556
rect 4897 6500 4953 6556
rect 4953 6500 4957 6556
rect 4893 6496 4957 6500
rect 4973 6556 5037 6560
rect 4973 6500 4977 6556
rect 4977 6500 5033 6556
rect 5033 6500 5037 6556
rect 4973 6496 5037 6500
rect 5053 6556 5117 6560
rect 5053 6500 5057 6556
rect 5057 6500 5113 6556
rect 5113 6500 5117 6556
rect 5053 6496 5117 6500
rect 6790 6556 6854 6560
rect 6790 6500 6794 6556
rect 6794 6500 6850 6556
rect 6850 6500 6854 6556
rect 6790 6496 6854 6500
rect 6870 6556 6934 6560
rect 6870 6500 6874 6556
rect 6874 6500 6930 6556
rect 6930 6500 6934 6556
rect 6870 6496 6934 6500
rect 6950 6556 7014 6560
rect 6950 6500 6954 6556
rect 6954 6500 7010 6556
rect 7010 6500 7014 6556
rect 6950 6496 7014 6500
rect 7030 6556 7094 6560
rect 7030 6500 7034 6556
rect 7034 6500 7090 6556
rect 7090 6500 7094 6556
rect 7030 6496 7094 6500
rect 8767 6556 8831 6560
rect 8767 6500 8771 6556
rect 8771 6500 8827 6556
rect 8827 6500 8831 6556
rect 8767 6496 8831 6500
rect 8847 6556 8911 6560
rect 8847 6500 8851 6556
rect 8851 6500 8907 6556
rect 8907 6500 8911 6556
rect 8847 6496 8911 6500
rect 8927 6556 8991 6560
rect 8927 6500 8931 6556
rect 8931 6500 8987 6556
rect 8987 6500 8991 6556
rect 8927 6496 8991 6500
rect 9007 6556 9071 6560
rect 9007 6500 9011 6556
rect 9011 6500 9067 6556
rect 9067 6500 9071 6556
rect 9007 6496 9071 6500
rect 1848 6012 1912 6016
rect 1848 5956 1852 6012
rect 1852 5956 1908 6012
rect 1908 5956 1912 6012
rect 1848 5952 1912 5956
rect 1928 6012 1992 6016
rect 1928 5956 1932 6012
rect 1932 5956 1988 6012
rect 1988 5956 1992 6012
rect 1928 5952 1992 5956
rect 2008 6012 2072 6016
rect 2008 5956 2012 6012
rect 2012 5956 2068 6012
rect 2068 5956 2072 6012
rect 2008 5952 2072 5956
rect 2088 6012 2152 6016
rect 2088 5956 2092 6012
rect 2092 5956 2148 6012
rect 2148 5956 2152 6012
rect 2088 5952 2152 5956
rect 3825 6012 3889 6016
rect 3825 5956 3829 6012
rect 3829 5956 3885 6012
rect 3885 5956 3889 6012
rect 3825 5952 3889 5956
rect 3905 6012 3969 6016
rect 3905 5956 3909 6012
rect 3909 5956 3965 6012
rect 3965 5956 3969 6012
rect 3905 5952 3969 5956
rect 3985 6012 4049 6016
rect 3985 5956 3989 6012
rect 3989 5956 4045 6012
rect 4045 5956 4049 6012
rect 3985 5952 4049 5956
rect 4065 6012 4129 6016
rect 4065 5956 4069 6012
rect 4069 5956 4125 6012
rect 4125 5956 4129 6012
rect 4065 5952 4129 5956
rect 5802 6012 5866 6016
rect 5802 5956 5806 6012
rect 5806 5956 5862 6012
rect 5862 5956 5866 6012
rect 5802 5952 5866 5956
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 7779 6012 7843 6016
rect 7779 5956 7783 6012
rect 7783 5956 7839 6012
rect 7839 5956 7843 6012
rect 7779 5952 7843 5956
rect 7859 6012 7923 6016
rect 7859 5956 7863 6012
rect 7863 5956 7919 6012
rect 7919 5956 7923 6012
rect 7859 5952 7923 5956
rect 7939 6012 8003 6016
rect 7939 5956 7943 6012
rect 7943 5956 7999 6012
rect 7999 5956 8003 6012
rect 7939 5952 8003 5956
rect 8019 6012 8083 6016
rect 8019 5956 8023 6012
rect 8023 5956 8079 6012
rect 8079 5956 8083 6012
rect 8019 5952 8083 5956
rect 2836 5468 2900 5472
rect 2836 5412 2840 5468
rect 2840 5412 2896 5468
rect 2896 5412 2900 5468
rect 2836 5408 2900 5412
rect 2916 5468 2980 5472
rect 2916 5412 2920 5468
rect 2920 5412 2976 5468
rect 2976 5412 2980 5468
rect 2916 5408 2980 5412
rect 2996 5468 3060 5472
rect 2996 5412 3000 5468
rect 3000 5412 3056 5468
rect 3056 5412 3060 5468
rect 2996 5408 3060 5412
rect 3076 5468 3140 5472
rect 3076 5412 3080 5468
rect 3080 5412 3136 5468
rect 3136 5412 3140 5468
rect 3076 5408 3140 5412
rect 4813 5468 4877 5472
rect 4813 5412 4817 5468
rect 4817 5412 4873 5468
rect 4873 5412 4877 5468
rect 4813 5408 4877 5412
rect 4893 5468 4957 5472
rect 4893 5412 4897 5468
rect 4897 5412 4953 5468
rect 4953 5412 4957 5468
rect 4893 5408 4957 5412
rect 4973 5468 5037 5472
rect 4973 5412 4977 5468
rect 4977 5412 5033 5468
rect 5033 5412 5037 5468
rect 4973 5408 5037 5412
rect 5053 5468 5117 5472
rect 5053 5412 5057 5468
rect 5057 5412 5113 5468
rect 5113 5412 5117 5468
rect 5053 5408 5117 5412
rect 6790 5468 6854 5472
rect 6790 5412 6794 5468
rect 6794 5412 6850 5468
rect 6850 5412 6854 5468
rect 6790 5408 6854 5412
rect 6870 5468 6934 5472
rect 6870 5412 6874 5468
rect 6874 5412 6930 5468
rect 6930 5412 6934 5468
rect 6870 5408 6934 5412
rect 6950 5468 7014 5472
rect 6950 5412 6954 5468
rect 6954 5412 7010 5468
rect 7010 5412 7014 5468
rect 6950 5408 7014 5412
rect 7030 5468 7094 5472
rect 7030 5412 7034 5468
rect 7034 5412 7090 5468
rect 7090 5412 7094 5468
rect 7030 5408 7094 5412
rect 8767 5468 8831 5472
rect 8767 5412 8771 5468
rect 8771 5412 8827 5468
rect 8827 5412 8831 5468
rect 8767 5408 8831 5412
rect 8847 5468 8911 5472
rect 8847 5412 8851 5468
rect 8851 5412 8907 5468
rect 8907 5412 8911 5468
rect 8847 5408 8911 5412
rect 8927 5468 8991 5472
rect 8927 5412 8931 5468
rect 8931 5412 8987 5468
rect 8987 5412 8991 5468
rect 8927 5408 8991 5412
rect 9007 5468 9071 5472
rect 9007 5412 9011 5468
rect 9011 5412 9067 5468
rect 9067 5412 9071 5468
rect 9007 5408 9071 5412
rect 1848 4924 1912 4928
rect 1848 4868 1852 4924
rect 1852 4868 1908 4924
rect 1908 4868 1912 4924
rect 1848 4864 1912 4868
rect 1928 4924 1992 4928
rect 1928 4868 1932 4924
rect 1932 4868 1988 4924
rect 1988 4868 1992 4924
rect 1928 4864 1992 4868
rect 2008 4924 2072 4928
rect 2008 4868 2012 4924
rect 2012 4868 2068 4924
rect 2068 4868 2072 4924
rect 2008 4864 2072 4868
rect 2088 4924 2152 4928
rect 2088 4868 2092 4924
rect 2092 4868 2148 4924
rect 2148 4868 2152 4924
rect 2088 4864 2152 4868
rect 3825 4924 3889 4928
rect 3825 4868 3829 4924
rect 3829 4868 3885 4924
rect 3885 4868 3889 4924
rect 3825 4864 3889 4868
rect 3905 4924 3969 4928
rect 3905 4868 3909 4924
rect 3909 4868 3965 4924
rect 3965 4868 3969 4924
rect 3905 4864 3969 4868
rect 3985 4924 4049 4928
rect 3985 4868 3989 4924
rect 3989 4868 4045 4924
rect 4045 4868 4049 4924
rect 3985 4864 4049 4868
rect 4065 4924 4129 4928
rect 4065 4868 4069 4924
rect 4069 4868 4125 4924
rect 4125 4868 4129 4924
rect 4065 4864 4129 4868
rect 5802 4924 5866 4928
rect 5802 4868 5806 4924
rect 5806 4868 5862 4924
rect 5862 4868 5866 4924
rect 5802 4864 5866 4868
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 7779 4924 7843 4928
rect 7779 4868 7783 4924
rect 7783 4868 7839 4924
rect 7839 4868 7843 4924
rect 7779 4864 7843 4868
rect 7859 4924 7923 4928
rect 7859 4868 7863 4924
rect 7863 4868 7919 4924
rect 7919 4868 7923 4924
rect 7859 4864 7923 4868
rect 7939 4924 8003 4928
rect 7939 4868 7943 4924
rect 7943 4868 7999 4924
rect 7999 4868 8003 4924
rect 7939 4864 8003 4868
rect 8019 4924 8083 4928
rect 8019 4868 8023 4924
rect 8023 4868 8079 4924
rect 8079 4868 8083 4924
rect 8019 4864 8083 4868
rect 2836 4380 2900 4384
rect 2836 4324 2840 4380
rect 2840 4324 2896 4380
rect 2896 4324 2900 4380
rect 2836 4320 2900 4324
rect 2916 4380 2980 4384
rect 2916 4324 2920 4380
rect 2920 4324 2976 4380
rect 2976 4324 2980 4380
rect 2916 4320 2980 4324
rect 2996 4380 3060 4384
rect 2996 4324 3000 4380
rect 3000 4324 3056 4380
rect 3056 4324 3060 4380
rect 2996 4320 3060 4324
rect 3076 4380 3140 4384
rect 3076 4324 3080 4380
rect 3080 4324 3136 4380
rect 3136 4324 3140 4380
rect 3076 4320 3140 4324
rect 4813 4380 4877 4384
rect 4813 4324 4817 4380
rect 4817 4324 4873 4380
rect 4873 4324 4877 4380
rect 4813 4320 4877 4324
rect 4893 4380 4957 4384
rect 4893 4324 4897 4380
rect 4897 4324 4953 4380
rect 4953 4324 4957 4380
rect 4893 4320 4957 4324
rect 4973 4380 5037 4384
rect 4973 4324 4977 4380
rect 4977 4324 5033 4380
rect 5033 4324 5037 4380
rect 4973 4320 5037 4324
rect 5053 4380 5117 4384
rect 5053 4324 5057 4380
rect 5057 4324 5113 4380
rect 5113 4324 5117 4380
rect 5053 4320 5117 4324
rect 6790 4380 6854 4384
rect 6790 4324 6794 4380
rect 6794 4324 6850 4380
rect 6850 4324 6854 4380
rect 6790 4320 6854 4324
rect 6870 4380 6934 4384
rect 6870 4324 6874 4380
rect 6874 4324 6930 4380
rect 6930 4324 6934 4380
rect 6870 4320 6934 4324
rect 6950 4380 7014 4384
rect 6950 4324 6954 4380
rect 6954 4324 7010 4380
rect 7010 4324 7014 4380
rect 6950 4320 7014 4324
rect 7030 4380 7094 4384
rect 7030 4324 7034 4380
rect 7034 4324 7090 4380
rect 7090 4324 7094 4380
rect 7030 4320 7094 4324
rect 8767 4380 8831 4384
rect 8767 4324 8771 4380
rect 8771 4324 8827 4380
rect 8827 4324 8831 4380
rect 8767 4320 8831 4324
rect 8847 4380 8911 4384
rect 8847 4324 8851 4380
rect 8851 4324 8907 4380
rect 8907 4324 8911 4380
rect 8847 4320 8911 4324
rect 8927 4380 8991 4384
rect 8927 4324 8931 4380
rect 8931 4324 8987 4380
rect 8987 4324 8991 4380
rect 8927 4320 8991 4324
rect 9007 4380 9071 4384
rect 9007 4324 9011 4380
rect 9011 4324 9067 4380
rect 9067 4324 9071 4380
rect 9007 4320 9071 4324
rect 1848 3836 1912 3840
rect 1848 3780 1852 3836
rect 1852 3780 1908 3836
rect 1908 3780 1912 3836
rect 1848 3776 1912 3780
rect 1928 3836 1992 3840
rect 1928 3780 1932 3836
rect 1932 3780 1988 3836
rect 1988 3780 1992 3836
rect 1928 3776 1992 3780
rect 2008 3836 2072 3840
rect 2008 3780 2012 3836
rect 2012 3780 2068 3836
rect 2068 3780 2072 3836
rect 2008 3776 2072 3780
rect 2088 3836 2152 3840
rect 2088 3780 2092 3836
rect 2092 3780 2148 3836
rect 2148 3780 2152 3836
rect 2088 3776 2152 3780
rect 3825 3836 3889 3840
rect 3825 3780 3829 3836
rect 3829 3780 3885 3836
rect 3885 3780 3889 3836
rect 3825 3776 3889 3780
rect 3905 3836 3969 3840
rect 3905 3780 3909 3836
rect 3909 3780 3965 3836
rect 3965 3780 3969 3836
rect 3905 3776 3969 3780
rect 3985 3836 4049 3840
rect 3985 3780 3989 3836
rect 3989 3780 4045 3836
rect 4045 3780 4049 3836
rect 3985 3776 4049 3780
rect 4065 3836 4129 3840
rect 4065 3780 4069 3836
rect 4069 3780 4125 3836
rect 4125 3780 4129 3836
rect 4065 3776 4129 3780
rect 5802 3836 5866 3840
rect 5802 3780 5806 3836
rect 5806 3780 5862 3836
rect 5862 3780 5866 3836
rect 5802 3776 5866 3780
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 7779 3836 7843 3840
rect 7779 3780 7783 3836
rect 7783 3780 7839 3836
rect 7839 3780 7843 3836
rect 7779 3776 7843 3780
rect 7859 3836 7923 3840
rect 7859 3780 7863 3836
rect 7863 3780 7919 3836
rect 7919 3780 7923 3836
rect 7859 3776 7923 3780
rect 7939 3836 8003 3840
rect 7939 3780 7943 3836
rect 7943 3780 7999 3836
rect 7999 3780 8003 3836
rect 7939 3776 8003 3780
rect 8019 3836 8083 3840
rect 8019 3780 8023 3836
rect 8023 3780 8079 3836
rect 8079 3780 8083 3836
rect 8019 3776 8083 3780
rect 2836 3292 2900 3296
rect 2836 3236 2840 3292
rect 2840 3236 2896 3292
rect 2896 3236 2900 3292
rect 2836 3232 2900 3236
rect 2916 3292 2980 3296
rect 2916 3236 2920 3292
rect 2920 3236 2976 3292
rect 2976 3236 2980 3292
rect 2916 3232 2980 3236
rect 2996 3292 3060 3296
rect 2996 3236 3000 3292
rect 3000 3236 3056 3292
rect 3056 3236 3060 3292
rect 2996 3232 3060 3236
rect 3076 3292 3140 3296
rect 3076 3236 3080 3292
rect 3080 3236 3136 3292
rect 3136 3236 3140 3292
rect 3076 3232 3140 3236
rect 4813 3292 4877 3296
rect 4813 3236 4817 3292
rect 4817 3236 4873 3292
rect 4873 3236 4877 3292
rect 4813 3232 4877 3236
rect 4893 3292 4957 3296
rect 4893 3236 4897 3292
rect 4897 3236 4953 3292
rect 4953 3236 4957 3292
rect 4893 3232 4957 3236
rect 4973 3292 5037 3296
rect 4973 3236 4977 3292
rect 4977 3236 5033 3292
rect 5033 3236 5037 3292
rect 4973 3232 5037 3236
rect 5053 3292 5117 3296
rect 5053 3236 5057 3292
rect 5057 3236 5113 3292
rect 5113 3236 5117 3292
rect 5053 3232 5117 3236
rect 6790 3292 6854 3296
rect 6790 3236 6794 3292
rect 6794 3236 6850 3292
rect 6850 3236 6854 3292
rect 6790 3232 6854 3236
rect 6870 3292 6934 3296
rect 6870 3236 6874 3292
rect 6874 3236 6930 3292
rect 6930 3236 6934 3292
rect 6870 3232 6934 3236
rect 6950 3292 7014 3296
rect 6950 3236 6954 3292
rect 6954 3236 7010 3292
rect 7010 3236 7014 3292
rect 6950 3232 7014 3236
rect 7030 3292 7094 3296
rect 7030 3236 7034 3292
rect 7034 3236 7090 3292
rect 7090 3236 7094 3292
rect 7030 3232 7094 3236
rect 8767 3292 8831 3296
rect 8767 3236 8771 3292
rect 8771 3236 8827 3292
rect 8827 3236 8831 3292
rect 8767 3232 8831 3236
rect 8847 3292 8911 3296
rect 8847 3236 8851 3292
rect 8851 3236 8907 3292
rect 8907 3236 8911 3292
rect 8847 3232 8911 3236
rect 8927 3292 8991 3296
rect 8927 3236 8931 3292
rect 8931 3236 8987 3292
rect 8987 3236 8991 3292
rect 8927 3232 8991 3236
rect 9007 3292 9071 3296
rect 9007 3236 9011 3292
rect 9011 3236 9067 3292
rect 9067 3236 9071 3292
rect 9007 3232 9071 3236
rect 1848 2748 1912 2752
rect 1848 2692 1852 2748
rect 1852 2692 1908 2748
rect 1908 2692 1912 2748
rect 1848 2688 1912 2692
rect 1928 2748 1992 2752
rect 1928 2692 1932 2748
rect 1932 2692 1988 2748
rect 1988 2692 1992 2748
rect 1928 2688 1992 2692
rect 2008 2748 2072 2752
rect 2008 2692 2012 2748
rect 2012 2692 2068 2748
rect 2068 2692 2072 2748
rect 2008 2688 2072 2692
rect 2088 2748 2152 2752
rect 2088 2692 2092 2748
rect 2092 2692 2148 2748
rect 2148 2692 2152 2748
rect 2088 2688 2152 2692
rect 3825 2748 3889 2752
rect 3825 2692 3829 2748
rect 3829 2692 3885 2748
rect 3885 2692 3889 2748
rect 3825 2688 3889 2692
rect 3905 2748 3969 2752
rect 3905 2692 3909 2748
rect 3909 2692 3965 2748
rect 3965 2692 3969 2748
rect 3905 2688 3969 2692
rect 3985 2748 4049 2752
rect 3985 2692 3989 2748
rect 3989 2692 4045 2748
rect 4045 2692 4049 2748
rect 3985 2688 4049 2692
rect 4065 2748 4129 2752
rect 4065 2692 4069 2748
rect 4069 2692 4125 2748
rect 4125 2692 4129 2748
rect 4065 2688 4129 2692
rect 5802 2748 5866 2752
rect 5802 2692 5806 2748
rect 5806 2692 5862 2748
rect 5862 2692 5866 2748
rect 5802 2688 5866 2692
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 7779 2748 7843 2752
rect 7779 2692 7783 2748
rect 7783 2692 7839 2748
rect 7839 2692 7843 2748
rect 7779 2688 7843 2692
rect 7859 2748 7923 2752
rect 7859 2692 7863 2748
rect 7863 2692 7919 2748
rect 7919 2692 7923 2748
rect 7859 2688 7923 2692
rect 7939 2748 8003 2752
rect 7939 2692 7943 2748
rect 7943 2692 7999 2748
rect 7999 2692 8003 2748
rect 7939 2688 8003 2692
rect 8019 2748 8083 2752
rect 8019 2692 8023 2748
rect 8023 2692 8079 2748
rect 8079 2692 8083 2748
rect 8019 2688 8083 2692
rect 2836 2204 2900 2208
rect 2836 2148 2840 2204
rect 2840 2148 2896 2204
rect 2896 2148 2900 2204
rect 2836 2144 2900 2148
rect 2916 2204 2980 2208
rect 2916 2148 2920 2204
rect 2920 2148 2976 2204
rect 2976 2148 2980 2204
rect 2916 2144 2980 2148
rect 2996 2204 3060 2208
rect 2996 2148 3000 2204
rect 3000 2148 3056 2204
rect 3056 2148 3060 2204
rect 2996 2144 3060 2148
rect 3076 2204 3140 2208
rect 3076 2148 3080 2204
rect 3080 2148 3136 2204
rect 3136 2148 3140 2204
rect 3076 2144 3140 2148
rect 4813 2204 4877 2208
rect 4813 2148 4817 2204
rect 4817 2148 4873 2204
rect 4873 2148 4877 2204
rect 4813 2144 4877 2148
rect 4893 2204 4957 2208
rect 4893 2148 4897 2204
rect 4897 2148 4953 2204
rect 4953 2148 4957 2204
rect 4893 2144 4957 2148
rect 4973 2204 5037 2208
rect 4973 2148 4977 2204
rect 4977 2148 5033 2204
rect 5033 2148 5037 2204
rect 4973 2144 5037 2148
rect 5053 2204 5117 2208
rect 5053 2148 5057 2204
rect 5057 2148 5113 2204
rect 5113 2148 5117 2204
rect 5053 2144 5117 2148
rect 6790 2204 6854 2208
rect 6790 2148 6794 2204
rect 6794 2148 6850 2204
rect 6850 2148 6854 2204
rect 6790 2144 6854 2148
rect 6870 2204 6934 2208
rect 6870 2148 6874 2204
rect 6874 2148 6930 2204
rect 6930 2148 6934 2204
rect 6870 2144 6934 2148
rect 6950 2204 7014 2208
rect 6950 2148 6954 2204
rect 6954 2148 7010 2204
rect 7010 2148 7014 2204
rect 6950 2144 7014 2148
rect 7030 2204 7094 2208
rect 7030 2148 7034 2204
rect 7034 2148 7090 2204
rect 7090 2148 7094 2204
rect 7030 2144 7094 2148
rect 8767 2204 8831 2208
rect 8767 2148 8771 2204
rect 8771 2148 8827 2204
rect 8827 2148 8831 2204
rect 8767 2144 8831 2148
rect 8847 2204 8911 2208
rect 8847 2148 8851 2204
rect 8851 2148 8907 2204
rect 8907 2148 8911 2204
rect 8847 2144 8911 2148
rect 8927 2204 8991 2208
rect 8927 2148 8931 2204
rect 8931 2148 8987 2204
rect 8987 2148 8991 2204
rect 8927 2144 8991 2148
rect 9007 2204 9071 2208
rect 9007 2148 9011 2204
rect 9011 2148 9067 2204
rect 9067 2148 9071 2204
rect 9007 2144 9071 2148
rect 1848 1660 1912 1664
rect 1848 1604 1852 1660
rect 1852 1604 1908 1660
rect 1908 1604 1912 1660
rect 1848 1600 1912 1604
rect 1928 1660 1992 1664
rect 1928 1604 1932 1660
rect 1932 1604 1988 1660
rect 1988 1604 1992 1660
rect 1928 1600 1992 1604
rect 2008 1660 2072 1664
rect 2008 1604 2012 1660
rect 2012 1604 2068 1660
rect 2068 1604 2072 1660
rect 2008 1600 2072 1604
rect 2088 1660 2152 1664
rect 2088 1604 2092 1660
rect 2092 1604 2148 1660
rect 2148 1604 2152 1660
rect 2088 1600 2152 1604
rect 3825 1660 3889 1664
rect 3825 1604 3829 1660
rect 3829 1604 3885 1660
rect 3885 1604 3889 1660
rect 3825 1600 3889 1604
rect 3905 1660 3969 1664
rect 3905 1604 3909 1660
rect 3909 1604 3965 1660
rect 3965 1604 3969 1660
rect 3905 1600 3969 1604
rect 3985 1660 4049 1664
rect 3985 1604 3989 1660
rect 3989 1604 4045 1660
rect 4045 1604 4049 1660
rect 3985 1600 4049 1604
rect 4065 1660 4129 1664
rect 4065 1604 4069 1660
rect 4069 1604 4125 1660
rect 4125 1604 4129 1660
rect 4065 1600 4129 1604
rect 5802 1660 5866 1664
rect 5802 1604 5806 1660
rect 5806 1604 5862 1660
rect 5862 1604 5866 1660
rect 5802 1600 5866 1604
rect 5882 1660 5946 1664
rect 5882 1604 5886 1660
rect 5886 1604 5942 1660
rect 5942 1604 5946 1660
rect 5882 1600 5946 1604
rect 5962 1660 6026 1664
rect 5962 1604 5966 1660
rect 5966 1604 6022 1660
rect 6022 1604 6026 1660
rect 5962 1600 6026 1604
rect 6042 1660 6106 1664
rect 6042 1604 6046 1660
rect 6046 1604 6102 1660
rect 6102 1604 6106 1660
rect 6042 1600 6106 1604
rect 7779 1660 7843 1664
rect 7779 1604 7783 1660
rect 7783 1604 7839 1660
rect 7839 1604 7843 1660
rect 7779 1600 7843 1604
rect 7859 1660 7923 1664
rect 7859 1604 7863 1660
rect 7863 1604 7919 1660
rect 7919 1604 7923 1660
rect 7859 1600 7923 1604
rect 7939 1660 8003 1664
rect 7939 1604 7943 1660
rect 7943 1604 7999 1660
rect 7999 1604 8003 1660
rect 7939 1600 8003 1604
rect 8019 1660 8083 1664
rect 8019 1604 8023 1660
rect 8023 1604 8079 1660
rect 8079 1604 8083 1660
rect 8019 1600 8083 1604
rect 2836 1116 2900 1120
rect 2836 1060 2840 1116
rect 2840 1060 2896 1116
rect 2896 1060 2900 1116
rect 2836 1056 2900 1060
rect 2916 1116 2980 1120
rect 2916 1060 2920 1116
rect 2920 1060 2976 1116
rect 2976 1060 2980 1116
rect 2916 1056 2980 1060
rect 2996 1116 3060 1120
rect 2996 1060 3000 1116
rect 3000 1060 3056 1116
rect 3056 1060 3060 1116
rect 2996 1056 3060 1060
rect 3076 1116 3140 1120
rect 3076 1060 3080 1116
rect 3080 1060 3136 1116
rect 3136 1060 3140 1116
rect 3076 1056 3140 1060
rect 4813 1116 4877 1120
rect 4813 1060 4817 1116
rect 4817 1060 4873 1116
rect 4873 1060 4877 1116
rect 4813 1056 4877 1060
rect 4893 1116 4957 1120
rect 4893 1060 4897 1116
rect 4897 1060 4953 1116
rect 4953 1060 4957 1116
rect 4893 1056 4957 1060
rect 4973 1116 5037 1120
rect 4973 1060 4977 1116
rect 4977 1060 5033 1116
rect 5033 1060 5037 1116
rect 4973 1056 5037 1060
rect 5053 1116 5117 1120
rect 5053 1060 5057 1116
rect 5057 1060 5113 1116
rect 5113 1060 5117 1116
rect 5053 1056 5117 1060
rect 6790 1116 6854 1120
rect 6790 1060 6794 1116
rect 6794 1060 6850 1116
rect 6850 1060 6854 1116
rect 6790 1056 6854 1060
rect 6870 1116 6934 1120
rect 6870 1060 6874 1116
rect 6874 1060 6930 1116
rect 6930 1060 6934 1116
rect 6870 1056 6934 1060
rect 6950 1116 7014 1120
rect 6950 1060 6954 1116
rect 6954 1060 7010 1116
rect 7010 1060 7014 1116
rect 6950 1056 7014 1060
rect 7030 1116 7094 1120
rect 7030 1060 7034 1116
rect 7034 1060 7090 1116
rect 7090 1060 7094 1116
rect 7030 1056 7094 1060
rect 8767 1116 8831 1120
rect 8767 1060 8771 1116
rect 8771 1060 8827 1116
rect 8827 1060 8831 1116
rect 8767 1056 8831 1060
rect 8847 1116 8911 1120
rect 8847 1060 8851 1116
rect 8851 1060 8907 1116
rect 8907 1060 8911 1116
rect 8847 1056 8911 1060
rect 8927 1116 8991 1120
rect 8927 1060 8931 1116
rect 8931 1060 8987 1116
rect 8987 1060 8991 1116
rect 8927 1056 8991 1060
rect 9007 1116 9071 1120
rect 9007 1060 9011 1116
rect 9011 1060 9067 1116
rect 9067 1060 9071 1116
rect 9007 1056 9071 1060
<< metal4 >>
rect 1840 14720 2160 14736
rect 1840 14656 1848 14720
rect 1912 14656 1928 14720
rect 1992 14656 2008 14720
rect 2072 14656 2088 14720
rect 2152 14656 2160 14720
rect 1840 13632 2160 14656
rect 1840 13568 1848 13632
rect 1912 13568 1928 13632
rect 1992 13568 2008 13632
rect 2072 13568 2088 13632
rect 2152 13568 2160 13632
rect 1840 12544 2160 13568
rect 1840 12480 1848 12544
rect 1912 12480 1928 12544
rect 1992 12480 2008 12544
rect 2072 12480 2088 12544
rect 2152 12480 2160 12544
rect 1840 11456 2160 12480
rect 1840 11392 1848 11456
rect 1912 11392 1928 11456
rect 1992 11392 2008 11456
rect 2072 11392 2088 11456
rect 2152 11392 2160 11456
rect 1840 10368 2160 11392
rect 1840 10304 1848 10368
rect 1912 10304 1928 10368
rect 1992 10304 2008 10368
rect 2072 10304 2088 10368
rect 2152 10304 2160 10368
rect 1840 9280 2160 10304
rect 1840 9216 1848 9280
rect 1912 9216 1928 9280
rect 1992 9216 2008 9280
rect 2072 9216 2088 9280
rect 2152 9216 2160 9280
rect 1840 8192 2160 9216
rect 1840 8128 1848 8192
rect 1912 8128 1928 8192
rect 1992 8128 2008 8192
rect 2072 8128 2088 8192
rect 2152 8128 2160 8192
rect 1840 7104 2160 8128
rect 1840 7040 1848 7104
rect 1912 7040 1928 7104
rect 1992 7040 2008 7104
rect 2072 7040 2088 7104
rect 2152 7040 2160 7104
rect 1840 6016 2160 7040
rect 1840 5952 1848 6016
rect 1912 5952 1928 6016
rect 1992 5952 2008 6016
rect 2072 5952 2088 6016
rect 2152 5952 2160 6016
rect 1840 4928 2160 5952
rect 1840 4864 1848 4928
rect 1912 4864 1928 4928
rect 1992 4864 2008 4928
rect 2072 4864 2088 4928
rect 2152 4864 2160 4928
rect 1840 3840 2160 4864
rect 1840 3776 1848 3840
rect 1912 3776 1928 3840
rect 1992 3776 2008 3840
rect 2072 3776 2088 3840
rect 2152 3776 2160 3840
rect 1840 2752 2160 3776
rect 1840 2688 1848 2752
rect 1912 2688 1928 2752
rect 1992 2688 2008 2752
rect 2072 2688 2088 2752
rect 2152 2688 2160 2752
rect 1840 1664 2160 2688
rect 1840 1600 1848 1664
rect 1912 1600 1928 1664
rect 1992 1600 2008 1664
rect 2072 1600 2088 1664
rect 2152 1600 2160 1664
rect 1840 1040 2160 1600
rect 2828 14176 3148 14736
rect 2828 14112 2836 14176
rect 2900 14112 2916 14176
rect 2980 14112 2996 14176
rect 3060 14112 3076 14176
rect 3140 14112 3148 14176
rect 2828 13088 3148 14112
rect 2828 13024 2836 13088
rect 2900 13024 2916 13088
rect 2980 13024 2996 13088
rect 3060 13024 3076 13088
rect 3140 13024 3148 13088
rect 2828 12000 3148 13024
rect 2828 11936 2836 12000
rect 2900 11936 2916 12000
rect 2980 11936 2996 12000
rect 3060 11936 3076 12000
rect 3140 11936 3148 12000
rect 2828 10912 3148 11936
rect 2828 10848 2836 10912
rect 2900 10848 2916 10912
rect 2980 10848 2996 10912
rect 3060 10848 3076 10912
rect 3140 10848 3148 10912
rect 2828 9824 3148 10848
rect 2828 9760 2836 9824
rect 2900 9760 2916 9824
rect 2980 9760 2996 9824
rect 3060 9760 3076 9824
rect 3140 9760 3148 9824
rect 2828 8736 3148 9760
rect 2828 8672 2836 8736
rect 2900 8672 2916 8736
rect 2980 8672 2996 8736
rect 3060 8672 3076 8736
rect 3140 8672 3148 8736
rect 2828 7648 3148 8672
rect 2828 7584 2836 7648
rect 2900 7584 2916 7648
rect 2980 7584 2996 7648
rect 3060 7584 3076 7648
rect 3140 7584 3148 7648
rect 2828 6560 3148 7584
rect 2828 6496 2836 6560
rect 2900 6496 2916 6560
rect 2980 6496 2996 6560
rect 3060 6496 3076 6560
rect 3140 6496 3148 6560
rect 2828 5472 3148 6496
rect 2828 5408 2836 5472
rect 2900 5408 2916 5472
rect 2980 5408 2996 5472
rect 3060 5408 3076 5472
rect 3140 5408 3148 5472
rect 2828 4384 3148 5408
rect 2828 4320 2836 4384
rect 2900 4320 2916 4384
rect 2980 4320 2996 4384
rect 3060 4320 3076 4384
rect 3140 4320 3148 4384
rect 2828 3296 3148 4320
rect 2828 3232 2836 3296
rect 2900 3232 2916 3296
rect 2980 3232 2996 3296
rect 3060 3232 3076 3296
rect 3140 3232 3148 3296
rect 2828 2208 3148 3232
rect 2828 2144 2836 2208
rect 2900 2144 2916 2208
rect 2980 2144 2996 2208
rect 3060 2144 3076 2208
rect 3140 2144 3148 2208
rect 2828 1120 3148 2144
rect 2828 1056 2836 1120
rect 2900 1056 2916 1120
rect 2980 1056 2996 1120
rect 3060 1056 3076 1120
rect 3140 1056 3148 1120
rect 2828 1040 3148 1056
rect 3817 14720 4137 14736
rect 3817 14656 3825 14720
rect 3889 14656 3905 14720
rect 3969 14656 3985 14720
rect 4049 14656 4065 14720
rect 4129 14656 4137 14720
rect 3817 13632 4137 14656
rect 3817 13568 3825 13632
rect 3889 13568 3905 13632
rect 3969 13568 3985 13632
rect 4049 13568 4065 13632
rect 4129 13568 4137 13632
rect 3817 12544 4137 13568
rect 3817 12480 3825 12544
rect 3889 12480 3905 12544
rect 3969 12480 3985 12544
rect 4049 12480 4065 12544
rect 4129 12480 4137 12544
rect 3817 11456 4137 12480
rect 3817 11392 3825 11456
rect 3889 11392 3905 11456
rect 3969 11392 3985 11456
rect 4049 11392 4065 11456
rect 4129 11392 4137 11456
rect 3817 10368 4137 11392
rect 3817 10304 3825 10368
rect 3889 10304 3905 10368
rect 3969 10304 3985 10368
rect 4049 10304 4065 10368
rect 4129 10304 4137 10368
rect 3817 9280 4137 10304
rect 3817 9216 3825 9280
rect 3889 9216 3905 9280
rect 3969 9216 3985 9280
rect 4049 9216 4065 9280
rect 4129 9216 4137 9280
rect 3817 8192 4137 9216
rect 3817 8128 3825 8192
rect 3889 8128 3905 8192
rect 3969 8128 3985 8192
rect 4049 8128 4065 8192
rect 4129 8128 4137 8192
rect 3817 7104 4137 8128
rect 3817 7040 3825 7104
rect 3889 7040 3905 7104
rect 3969 7040 3985 7104
rect 4049 7040 4065 7104
rect 4129 7040 4137 7104
rect 3817 6016 4137 7040
rect 3817 5952 3825 6016
rect 3889 5952 3905 6016
rect 3969 5952 3985 6016
rect 4049 5952 4065 6016
rect 4129 5952 4137 6016
rect 3817 4928 4137 5952
rect 3817 4864 3825 4928
rect 3889 4864 3905 4928
rect 3969 4864 3985 4928
rect 4049 4864 4065 4928
rect 4129 4864 4137 4928
rect 3817 3840 4137 4864
rect 3817 3776 3825 3840
rect 3889 3776 3905 3840
rect 3969 3776 3985 3840
rect 4049 3776 4065 3840
rect 4129 3776 4137 3840
rect 3817 2752 4137 3776
rect 3817 2688 3825 2752
rect 3889 2688 3905 2752
rect 3969 2688 3985 2752
rect 4049 2688 4065 2752
rect 4129 2688 4137 2752
rect 3817 1664 4137 2688
rect 3817 1600 3825 1664
rect 3889 1600 3905 1664
rect 3969 1600 3985 1664
rect 4049 1600 4065 1664
rect 4129 1600 4137 1664
rect 3817 1040 4137 1600
rect 4805 14176 5125 14736
rect 4805 14112 4813 14176
rect 4877 14112 4893 14176
rect 4957 14112 4973 14176
rect 5037 14112 5053 14176
rect 5117 14112 5125 14176
rect 4805 13088 5125 14112
rect 4805 13024 4813 13088
rect 4877 13024 4893 13088
rect 4957 13024 4973 13088
rect 5037 13024 5053 13088
rect 5117 13024 5125 13088
rect 4805 12000 5125 13024
rect 4805 11936 4813 12000
rect 4877 11936 4893 12000
rect 4957 11936 4973 12000
rect 5037 11936 5053 12000
rect 5117 11936 5125 12000
rect 4805 10912 5125 11936
rect 4805 10848 4813 10912
rect 4877 10848 4893 10912
rect 4957 10848 4973 10912
rect 5037 10848 5053 10912
rect 5117 10848 5125 10912
rect 4805 9824 5125 10848
rect 4805 9760 4813 9824
rect 4877 9760 4893 9824
rect 4957 9760 4973 9824
rect 5037 9760 5053 9824
rect 5117 9760 5125 9824
rect 4805 8736 5125 9760
rect 4805 8672 4813 8736
rect 4877 8672 4893 8736
rect 4957 8672 4973 8736
rect 5037 8672 5053 8736
rect 5117 8672 5125 8736
rect 4805 7648 5125 8672
rect 4805 7584 4813 7648
rect 4877 7584 4893 7648
rect 4957 7584 4973 7648
rect 5037 7584 5053 7648
rect 5117 7584 5125 7648
rect 4805 6560 5125 7584
rect 4805 6496 4813 6560
rect 4877 6496 4893 6560
rect 4957 6496 4973 6560
rect 5037 6496 5053 6560
rect 5117 6496 5125 6560
rect 4805 5472 5125 6496
rect 4805 5408 4813 5472
rect 4877 5408 4893 5472
rect 4957 5408 4973 5472
rect 5037 5408 5053 5472
rect 5117 5408 5125 5472
rect 4805 4384 5125 5408
rect 4805 4320 4813 4384
rect 4877 4320 4893 4384
rect 4957 4320 4973 4384
rect 5037 4320 5053 4384
rect 5117 4320 5125 4384
rect 4805 3296 5125 4320
rect 4805 3232 4813 3296
rect 4877 3232 4893 3296
rect 4957 3232 4973 3296
rect 5037 3232 5053 3296
rect 5117 3232 5125 3296
rect 4805 2208 5125 3232
rect 4805 2144 4813 2208
rect 4877 2144 4893 2208
rect 4957 2144 4973 2208
rect 5037 2144 5053 2208
rect 5117 2144 5125 2208
rect 4805 1120 5125 2144
rect 4805 1056 4813 1120
rect 4877 1056 4893 1120
rect 4957 1056 4973 1120
rect 5037 1056 5053 1120
rect 5117 1056 5125 1120
rect 4805 1040 5125 1056
rect 5794 14720 6114 14736
rect 5794 14656 5802 14720
rect 5866 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6114 14720
rect 5794 13632 6114 14656
rect 5794 13568 5802 13632
rect 5866 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6114 13632
rect 5794 12544 6114 13568
rect 5794 12480 5802 12544
rect 5866 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6114 12544
rect 5794 11456 6114 12480
rect 5794 11392 5802 11456
rect 5866 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6114 11456
rect 5794 10368 6114 11392
rect 5794 10304 5802 10368
rect 5866 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6114 10368
rect 5794 9280 6114 10304
rect 5794 9216 5802 9280
rect 5866 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6114 9280
rect 5794 8192 6114 9216
rect 5794 8128 5802 8192
rect 5866 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6114 8192
rect 5794 7104 6114 8128
rect 5794 7040 5802 7104
rect 5866 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6114 7104
rect 5794 6016 6114 7040
rect 5794 5952 5802 6016
rect 5866 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6114 6016
rect 5794 4928 6114 5952
rect 5794 4864 5802 4928
rect 5866 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6114 4928
rect 5794 3840 6114 4864
rect 5794 3776 5802 3840
rect 5866 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6114 3840
rect 5794 2752 6114 3776
rect 5794 2688 5802 2752
rect 5866 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6114 2752
rect 5794 1664 6114 2688
rect 5794 1600 5802 1664
rect 5866 1600 5882 1664
rect 5946 1600 5962 1664
rect 6026 1600 6042 1664
rect 6106 1600 6114 1664
rect 5794 1040 6114 1600
rect 6782 14176 7102 14736
rect 6782 14112 6790 14176
rect 6854 14112 6870 14176
rect 6934 14112 6950 14176
rect 7014 14112 7030 14176
rect 7094 14112 7102 14176
rect 6782 13088 7102 14112
rect 6782 13024 6790 13088
rect 6854 13024 6870 13088
rect 6934 13024 6950 13088
rect 7014 13024 7030 13088
rect 7094 13024 7102 13088
rect 6782 12000 7102 13024
rect 6782 11936 6790 12000
rect 6854 11936 6870 12000
rect 6934 11936 6950 12000
rect 7014 11936 7030 12000
rect 7094 11936 7102 12000
rect 6782 10912 7102 11936
rect 6782 10848 6790 10912
rect 6854 10848 6870 10912
rect 6934 10848 6950 10912
rect 7014 10848 7030 10912
rect 7094 10848 7102 10912
rect 6782 9824 7102 10848
rect 6782 9760 6790 9824
rect 6854 9760 6870 9824
rect 6934 9760 6950 9824
rect 7014 9760 7030 9824
rect 7094 9760 7102 9824
rect 6782 8736 7102 9760
rect 6782 8672 6790 8736
rect 6854 8672 6870 8736
rect 6934 8672 6950 8736
rect 7014 8672 7030 8736
rect 7094 8672 7102 8736
rect 6782 7648 7102 8672
rect 6782 7584 6790 7648
rect 6854 7584 6870 7648
rect 6934 7584 6950 7648
rect 7014 7584 7030 7648
rect 7094 7584 7102 7648
rect 6782 6560 7102 7584
rect 6782 6496 6790 6560
rect 6854 6496 6870 6560
rect 6934 6496 6950 6560
rect 7014 6496 7030 6560
rect 7094 6496 7102 6560
rect 6782 5472 7102 6496
rect 6782 5408 6790 5472
rect 6854 5408 6870 5472
rect 6934 5408 6950 5472
rect 7014 5408 7030 5472
rect 7094 5408 7102 5472
rect 6782 4384 7102 5408
rect 6782 4320 6790 4384
rect 6854 4320 6870 4384
rect 6934 4320 6950 4384
rect 7014 4320 7030 4384
rect 7094 4320 7102 4384
rect 6782 3296 7102 4320
rect 6782 3232 6790 3296
rect 6854 3232 6870 3296
rect 6934 3232 6950 3296
rect 7014 3232 7030 3296
rect 7094 3232 7102 3296
rect 6782 2208 7102 3232
rect 6782 2144 6790 2208
rect 6854 2144 6870 2208
rect 6934 2144 6950 2208
rect 7014 2144 7030 2208
rect 7094 2144 7102 2208
rect 6782 1120 7102 2144
rect 6782 1056 6790 1120
rect 6854 1056 6870 1120
rect 6934 1056 6950 1120
rect 7014 1056 7030 1120
rect 7094 1056 7102 1120
rect 6782 1040 7102 1056
rect 7771 14720 8091 14736
rect 7771 14656 7779 14720
rect 7843 14656 7859 14720
rect 7923 14656 7939 14720
rect 8003 14656 8019 14720
rect 8083 14656 8091 14720
rect 7771 13632 8091 14656
rect 7771 13568 7779 13632
rect 7843 13568 7859 13632
rect 7923 13568 7939 13632
rect 8003 13568 8019 13632
rect 8083 13568 8091 13632
rect 7771 12544 8091 13568
rect 7771 12480 7779 12544
rect 7843 12480 7859 12544
rect 7923 12480 7939 12544
rect 8003 12480 8019 12544
rect 8083 12480 8091 12544
rect 7771 11456 8091 12480
rect 7771 11392 7779 11456
rect 7843 11392 7859 11456
rect 7923 11392 7939 11456
rect 8003 11392 8019 11456
rect 8083 11392 8091 11456
rect 7771 10368 8091 11392
rect 7771 10304 7779 10368
rect 7843 10304 7859 10368
rect 7923 10304 7939 10368
rect 8003 10304 8019 10368
rect 8083 10304 8091 10368
rect 7771 9280 8091 10304
rect 7771 9216 7779 9280
rect 7843 9216 7859 9280
rect 7923 9216 7939 9280
rect 8003 9216 8019 9280
rect 8083 9216 8091 9280
rect 7771 8192 8091 9216
rect 7771 8128 7779 8192
rect 7843 8128 7859 8192
rect 7923 8128 7939 8192
rect 8003 8128 8019 8192
rect 8083 8128 8091 8192
rect 7771 7104 8091 8128
rect 7771 7040 7779 7104
rect 7843 7040 7859 7104
rect 7923 7040 7939 7104
rect 8003 7040 8019 7104
rect 8083 7040 8091 7104
rect 7771 6016 8091 7040
rect 7771 5952 7779 6016
rect 7843 5952 7859 6016
rect 7923 5952 7939 6016
rect 8003 5952 8019 6016
rect 8083 5952 8091 6016
rect 7771 4928 8091 5952
rect 7771 4864 7779 4928
rect 7843 4864 7859 4928
rect 7923 4864 7939 4928
rect 8003 4864 8019 4928
rect 8083 4864 8091 4928
rect 7771 3840 8091 4864
rect 7771 3776 7779 3840
rect 7843 3776 7859 3840
rect 7923 3776 7939 3840
rect 8003 3776 8019 3840
rect 8083 3776 8091 3840
rect 7771 2752 8091 3776
rect 7771 2688 7779 2752
rect 7843 2688 7859 2752
rect 7923 2688 7939 2752
rect 8003 2688 8019 2752
rect 8083 2688 8091 2752
rect 7771 1664 8091 2688
rect 7771 1600 7779 1664
rect 7843 1600 7859 1664
rect 7923 1600 7939 1664
rect 8003 1600 8019 1664
rect 8083 1600 8091 1664
rect 7771 1040 8091 1600
rect 8759 14176 9079 14736
rect 8759 14112 8767 14176
rect 8831 14112 8847 14176
rect 8911 14112 8927 14176
rect 8991 14112 9007 14176
rect 9071 14112 9079 14176
rect 8759 13088 9079 14112
rect 8759 13024 8767 13088
rect 8831 13024 8847 13088
rect 8911 13024 8927 13088
rect 8991 13024 9007 13088
rect 9071 13024 9079 13088
rect 8759 12000 9079 13024
rect 8759 11936 8767 12000
rect 8831 11936 8847 12000
rect 8911 11936 8927 12000
rect 8991 11936 9007 12000
rect 9071 11936 9079 12000
rect 8759 10912 9079 11936
rect 8759 10848 8767 10912
rect 8831 10848 8847 10912
rect 8911 10848 8927 10912
rect 8991 10848 9007 10912
rect 9071 10848 9079 10912
rect 8759 9824 9079 10848
rect 8759 9760 8767 9824
rect 8831 9760 8847 9824
rect 8911 9760 8927 9824
rect 8991 9760 9007 9824
rect 9071 9760 9079 9824
rect 8759 8736 9079 9760
rect 8759 8672 8767 8736
rect 8831 8672 8847 8736
rect 8911 8672 8927 8736
rect 8991 8672 9007 8736
rect 9071 8672 9079 8736
rect 8759 7648 9079 8672
rect 8759 7584 8767 7648
rect 8831 7584 8847 7648
rect 8911 7584 8927 7648
rect 8991 7584 9007 7648
rect 9071 7584 9079 7648
rect 8759 6560 9079 7584
rect 8759 6496 8767 6560
rect 8831 6496 8847 6560
rect 8911 6496 8927 6560
rect 8991 6496 9007 6560
rect 9071 6496 9079 6560
rect 8759 5472 9079 6496
rect 8759 5408 8767 5472
rect 8831 5408 8847 5472
rect 8911 5408 8927 5472
rect 8991 5408 9007 5472
rect 9071 5408 9079 5472
rect 8759 4384 9079 5408
rect 8759 4320 8767 4384
rect 8831 4320 8847 4384
rect 8911 4320 8927 4384
rect 8991 4320 9007 4384
rect 9071 4320 9079 4384
rect 8759 3296 9079 4320
rect 8759 3232 8767 3296
rect 8831 3232 8847 3296
rect 8911 3232 8927 3296
rect 8991 3232 9007 3296
rect 9071 3232 9079 3296
rect 8759 2208 9079 3232
rect 8759 2144 8767 2208
rect 8831 2144 8847 2208
rect 8911 2144 8927 2208
rect 8991 2144 9007 2208
rect 9071 2144 9079 2208
rect 8759 1120 9079 2144
rect 8759 1056 8767 1120
rect 8831 1056 8847 1120
rect 8911 1056 8927 1120
rect 8991 1056 9007 1120
rect 9071 1056 9079 1120
rect 8759 1040 9079 1056
use sky130_fd_sc_hd__nor2_4  _06_
timestamp 1750019440
transform 1 0 7820 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _07_
timestamp 1750019440
transform -1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1750019440
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _09_
timestamp 1750019440
transform -1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1750019440
transform -1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 1750019440
transform -1 0 8556 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1750019440
transform -1 0 8096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _13_
timestamp 1750019440
transform -1 0 8556 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1750019440
transform -1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _15_
timestamp 1750019440
transform -1 0 8556 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1750019440
transform -1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _17_
timestamp 1750019440
transform 1 0 8004 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1750019440
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _19_
timestamp 1750019440
transform -1 0 8648 0 -1 11968
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1750019440
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15
timestamp 1750019440
transform 1 0 2392 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_23
timestamp 1750019440
transform 1 0 3128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1750019440
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1750019440
transform 1 0 3680 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1750019440
transform 1 0 4784 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1750019440
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1750019440
transform 1 0 6256 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69
timestamp 1750019440
transform 1 0 7360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_75
timestamp 1750019440
transform 1 0 7912 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1750019440
transform 1 0 1288 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1750019440
transform 1 0 2392 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1750019440
transform 1 0 3496 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1750019440
transform 1 0 4600 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1750019440
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1750019440
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1750019440
transform 1 0 6256 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_69
timestamp 1750019440
transform 1 0 7360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 1750019440
transform 1 0 7728 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1750019440
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1750019440
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1750019440
transform 1 0 3496 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1750019440
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1750019440
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1750019440
transform 1 0 5888 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1750019440
transform 1 0 6992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1750019440
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1750019440
transform 1 0 1288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1750019440
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1750019440
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1750019440
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1750019440
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1750019440
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1750019440
transform 1 0 6256 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 1750019440
transform 1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_81
timestamp 1750019440
transform 1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1750019440
transform 1 0 1288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1750019440
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1750019440
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1750019440
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1750019440
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1750019440
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1750019440
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1750019440
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1750019440
transform 1 0 1288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1750019440
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1750019440
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1750019440
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1750019440
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1750019440
transform 1 0 6072 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1750019440
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1750019440
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_81
timestamp 1750019440
transform 1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1750019440
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1750019440
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1750019440
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1750019440
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1750019440
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1750019440
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1750019440
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1750019440
transform 1 0 8096 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1750019440
transform 1 0 1288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1750019440
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1750019440
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1750019440
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1750019440
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1750019440
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1750019440
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_69
timestamp 1750019440
transform 1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_82
timestamp 1750019440
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1750019440
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1750019440
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1750019440
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1750019440
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1750019440
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1750019440
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1750019440
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1750019440
transform 1 0 8096 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1750019440
transform 1 0 1288 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1750019440
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1750019440
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1750019440
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1750019440
transform 1 0 5704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1750019440
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1750019440
transform 1 0 6256 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1750019440
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_81
timestamp 1750019440
transform 1 0 8464 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1750019440
transform 1 0 1288 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1750019440
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1750019440
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1750019440
transform 1 0 3680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1750019440
transform 1 0 4784 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1750019440
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 1750019440
transform 1 0 6992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_82
timestamp 1750019440
transform 1 0 8556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1750019440
transform 1 0 1288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1750019440
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1750019440
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1750019440
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1750019440
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1750019440
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1750019440
transform 1 0 6256 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1750019440
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_81
timestamp 1750019440
transform 1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1750019440
transform 1 0 1288 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1750019440
transform 1 0 2392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1750019440
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1750019440
transform 1 0 3680 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1750019440
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1750019440
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1750019440
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1750019440
transform 1 0 8096 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1750019440
transform 1 0 1288 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1750019440
transform 1 0 2392 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1750019440
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1750019440
transform 1 0 4600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1750019440
transform 1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1750019440
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1750019440
transform 1 0 6256 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1750019440
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_81
timestamp 1750019440
transform 1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1750019440
transform 1 0 1288 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1750019440
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1750019440
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1750019440
transform 1 0 3680 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1750019440
transform 1 0 4784 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1750019440
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_65
timestamp 1750019440
transform 1 0 6992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_82
timestamp 1750019440
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1750019440
transform 1 0 1288 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1750019440
transform 1 0 2392 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1750019440
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1750019440
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1750019440
transform 1 0 5704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1750019440
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1750019440
transform 1 0 6256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1750019440
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_81
timestamp 1750019440
transform 1 0 8464 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1750019440
transform 1 0 1288 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1750019440
transform 1 0 2392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1750019440
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1750019440
transform 1 0 3680 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1750019440
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1750019440
transform 1 0 5888 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1750019440
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1750019440
transform 1 0 8096 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1750019440
transform 1 0 1288 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1750019440
transform 1 0 2392 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1750019440
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1750019440
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1750019440
transform 1 0 5704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1750019440
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1750019440
transform 1 0 6256 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_69
timestamp 1750019440
transform 1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_82
timestamp 1750019440
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1750019440
transform 1 0 1288 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1750019440
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1750019440
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1750019440
transform 1 0 3680 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1750019440
transform 1 0 4784 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1750019440
transform 1 0 5888 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp 1750019440
transform 1 0 6992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_73
timestamp 1750019440
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_82
timestamp 1750019440
transform 1 0 8556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1750019440
transform 1 0 1288 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1750019440
transform 1 0 2392 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1750019440
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1750019440
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1750019440
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1750019440
transform 1 0 6072 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1750019440
transform 1 0 6256 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_69
timestamp 1750019440
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_73
timestamp 1750019440
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1750019440
transform 1 0 1288 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1750019440
transform 1 0 2392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1750019440
transform 1 0 3496 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1750019440
transform 1 0 3680 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1750019440
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1750019440
transform 1 0 5888 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1750019440
transform 1 0 6992 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_77
timestamp 1750019440
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1750019440
transform 1 0 1288 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1750019440
transform 1 0 2392 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1750019440
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1750019440
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1750019440
transform 1 0 5704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1750019440
transform 1 0 6072 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1750019440
transform 1 0 6256 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1750019440
transform 1 0 7360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_81
timestamp 1750019440
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1750019440
transform 1 0 1288 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1750019440
transform 1 0 2392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1750019440
transform 1 0 3496 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1750019440
transform 1 0 3680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1750019440
transform 1 0 4784 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1750019440
transform 1 0 5888 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1750019440
transform 1 0 6992 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1750019440
transform 1 0 8096 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1750019440
transform 1 0 1288 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1750019440
transform 1 0 2392 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1750019440
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1750019440
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1750019440
transform 1 0 5704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1750019440
transform 1 0 6072 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1750019440
transform 1 0 6256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1750019440
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_81
timestamp 1750019440
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1750019440
transform 1 0 1288 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1750019440
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1750019440
transform 1 0 3496 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1750019440
transform 1 0 3680 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1750019440
transform 1 0 4784 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_53
timestamp 1750019440
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_57
timestamp 1750019440
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_69
timestamp 1750019440
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_81
timestamp 1750019440
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1749572018
transform 1 0 2576 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1750019440
transform 1 0 7544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_25
timestamp 1750019440
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1750019440
transform -1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_26
timestamp 1750019440
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1750019440
transform -1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_27
timestamp 1750019440
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1750019440
transform -1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_28
timestamp 1750019440
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1750019440
transform -1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_29
timestamp 1750019440
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1750019440
transform -1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_30
timestamp 1750019440
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1750019440
transform -1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_31
timestamp 1750019440
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1750019440
transform -1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_32
timestamp 1750019440
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1750019440
transform -1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_33
timestamp 1750019440
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1750019440
transform -1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_34
timestamp 1750019440
transform 1 0 1012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1750019440
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_35
timestamp 1750019440
transform 1 0 1012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1750019440
transform -1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_36
timestamp 1750019440
transform 1 0 1012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1750019440
transform -1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_37
timestamp 1750019440
transform 1 0 1012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1750019440
transform -1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_38
timestamp 1750019440
transform 1 0 1012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1750019440
transform -1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_39
timestamp 1750019440
transform 1 0 1012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1750019440
transform -1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_40
timestamp 1750019440
transform 1 0 1012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1750019440
transform -1 0 8924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_41
timestamp 1750019440
transform 1 0 1012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1750019440
transform -1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_42
timestamp 1750019440
transform 1 0 1012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1750019440
transform -1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_43
timestamp 1750019440
transform 1 0 1012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1750019440
transform -1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_44
timestamp 1750019440
transform 1 0 1012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1750019440
transform -1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_45
timestamp 1750019440
transform 1 0 1012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1750019440
transform -1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_46
timestamp 1750019440
transform 1 0 1012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1750019440
transform -1 0 8924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_47
timestamp 1750019440
transform 1 0 1012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1750019440
transform -1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_48
timestamp 1750019440
transform 1 0 1012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1750019440
transform -1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_49
timestamp 1750019440
transform 1 0 1012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1750019440
transform -1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp 1750019440
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp 1750019440
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_52
timestamp 1750019440
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 1750019440
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp 1750019440
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp 1750019440
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_56
timestamp 1750019440
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1750019440
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_58
timestamp 1750019440
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp 1750019440
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp 1750019440
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_61
timestamp 1750019440
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_62
timestamp 1750019440
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_63
timestamp 1750019440
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_64
timestamp 1750019440
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_65
timestamp 1750019440
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_66
timestamp 1750019440
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_67
timestamp 1750019440
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_68
timestamp 1750019440
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_69
timestamp 1750019440
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_70
timestamp 1750019440
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_71
timestamp 1750019440
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_72
timestamp 1750019440
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_73
timestamp 1750019440
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_74
timestamp 1750019440
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_75
timestamp 1750019440
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_76
timestamp 1750019440
transform 1 0 6164 0 1 14144
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5045 14144 5045 14144 4 VGND
rlabel metal1 s 4968 14688 4968 14688 4 VPWR
rlabel metal1 s 7912 3026 7912 3026 4 _00_
rlabel metal1 s 7958 5168 7958 5168 4 _01_
rlabel metal1 s 8096 6766 8096 6766 4 _02_
rlabel metal1 s 8096 8942 8096 8942 4 _03_
rlabel metal1 s 8004 10642 8004 10642 4 _04_
rlabel metal2 s 8510 11764 8510 11764 4 _05_
rlabel metal2 s 2530 806 2530 806 4 a
rlabel metal2 s 7498 840 7498 840 4 b
rlabel metal3 s 9484 1156 9484 1156 4 n[0]
rlabel metal2 s 7682 3111 7682 3111 4 n[1]
rlabel metal3 s 8932 4964 8932 4964 4 n[2]
rlabel metal2 s 7866 6749 7866 6749 4 n[3]
rlabel metal2 s 8326 1700 8326 1700 4 net1
rlabel metal1 s 8372 8942 8372 8942 4 net2
rlabel metal3 s 9461 8772 9461 8772 4 p[0]
rlabel metal2 s 7774 10727 7774 10727 4 p[1]
rlabel metal1 s 8372 12410 8372 12410 4 p[2]
rlabel metal1 s 8188 11730 8188 11730 4 p[3]
flabel metal4 s 8759 1040 9079 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6782 1040 7102 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4805 1040 5125 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2828 1040 3148 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7771 1040 8091 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5794 1040 6114 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3817 1040 4137 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1840 1040 2160 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 2502 0 2558 400 0 FreeSans 280 90 0 0 a
port 3 nsew
flabel metal2 s 7470 0 7526 400 0 FreeSans 280 90 0 0 b
port 4 nsew
flabel metal3 s 9600 1096 10000 1216 0 FreeSans 600 0 0 0 n[0]
port 5 nsew
flabel metal3 s 9600 3000 10000 3120 0 FreeSans 600 0 0 0 n[1]
port 6 nsew
flabel metal3 s 9600 4904 10000 5024 0 FreeSans 600 0 0 0 n[2]
port 7 nsew
flabel metal3 s 9600 6808 10000 6928 0 FreeSans 600 0 0 0 n[3]
port 8 nsew
flabel metal3 s 9600 8712 10000 8832 0 FreeSans 600 0 0 0 p[0]
port 9 nsew
flabel metal3 s 9600 10616 10000 10736 0 FreeSans 600 0 0 0 p[1]
port 10 nsew
flabel metal3 s 9600 12520 10000 12640 0 FreeSans 600 0 0 0 p[2]
port 11 nsew
flabel metal3 s 9600 14424 10000 14544 0 FreeSans 600 0 0 0 p[3]
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 16000
string GDS_END 219294
string GDS_FILE ../gds/Decoder.gds
string GDS_START 64426
<< end >>
