magic
tech sky130A
magscale 1 2
timestamp 1750689032
<< metal1 >>
rect 27670 43910 27726 43916
rect 19124 43775 19193 43781
rect 19193 43706 26029 43775
rect 26098 43706 26104 43775
rect 19124 43700 19193 43706
rect 27670 42902 27726 43854
rect 27664 42846 27670 42902
rect 27726 42846 27732 42902
rect 19227 41739 19293 41745
rect 27107 41739 27173 41745
rect 12793 41673 12799 41739
rect 12865 41673 19227 41739
rect 23387 41673 23393 41739
rect 23459 41673 27107 41739
rect 19227 41667 19293 41673
rect 27107 41667 27173 41673
rect 23618 40916 23674 40922
rect 10994 40844 11000 40900
rect 11056 40844 11062 40900
rect 19420 40860 19426 40916
rect 19482 40860 23618 40916
rect 23618 40854 23674 40860
rect 6026 40646 6032 40702
rect 6088 40646 6094 40702
rect 6032 38848 6088 40646
rect 11000 38954 11056 40844
rect 10994 38898 11000 38954
rect 11056 38898 11062 38954
rect 6032 38770 6088 38792
rect -32 -26 -26 26
rect 26 -26 32 26
<< via1 >>
rect 27670 43854 27726 43910
rect 19124 43706 19193 43775
rect 26029 43706 26098 43775
rect 27670 42846 27726 42902
rect 12799 41673 12865 41739
rect 19227 41673 19293 41739
rect 23393 41673 23459 41739
rect 27107 41673 27173 41739
rect 11000 40844 11056 40900
rect 19426 40860 19482 40916
rect 23618 40860 23674 40916
rect 6032 40646 6088 40702
rect 11000 38898 11056 38954
rect 6032 38792 6088 38848
rect -26 -26 26 26
<< metal2 >>
rect 28214 44406 28274 44408
rect 28207 44350 28216 44406
rect 28272 44350 28281 44406
rect 7238 44164 7298 44166
rect 7231 44108 7240 44164
rect 7296 44108 7305 44164
rect 6686 44082 6746 44084
rect 6679 44026 6688 44082
rect 6744 44026 6753 44082
rect 6130 43982 6199 43987
rect 6126 43923 6135 43982
rect 6194 43923 6203 43982
rect 6130 43775 6199 43923
rect 6686 43775 6746 44026
rect 7238 43775 7298 44108
rect 7790 44042 7850 44044
rect 7783 43986 7792 44042
rect 7848 43986 7857 44042
rect 18830 44024 18890 44026
rect 7790 43775 7850 43986
rect 16070 43976 16130 43978
rect 8894 43972 8954 43974
rect 8342 43962 8402 43964
rect 8335 43906 8344 43962
rect 8400 43906 8409 43962
rect 8887 43916 8896 43972
rect 8952 43916 8961 43972
rect 12758 43966 12818 43968
rect 10000 43958 10056 43965
rect 12206 43958 12266 43960
rect 9998 43956 10058 43958
rect 11654 43956 11714 43958
rect 9446 43940 9506 43942
rect 8342 43775 8402 43906
rect 8894 43775 8954 43916
rect 9439 43884 9448 43940
rect 9504 43884 9513 43940
rect 9998 43900 10000 43956
rect 10056 43900 10058 43956
rect 10550 43930 10610 43932
rect 9446 43775 9506 43884
rect 9998 43775 10058 43900
rect 10543 43874 10552 43930
rect 10608 43874 10617 43930
rect 11102 43904 11162 43906
rect 10550 43775 10610 43874
rect 11095 43848 11104 43904
rect 11160 43848 11169 43904
rect 11647 43900 11656 43956
rect 11712 43900 11721 43956
rect 12199 43902 12208 43958
rect 12264 43902 12273 43958
rect 12751 43910 12760 43966
rect 12816 43910 12825 43966
rect 13862 43950 13922 43952
rect 13310 43934 13370 43936
rect 11102 43775 11162 43848
rect 11654 43775 11714 43900
rect 12206 43775 12266 43902
rect 12758 43775 12818 43910
rect 13303 43878 13312 43934
rect 13368 43878 13377 43934
rect 13855 43894 13864 43950
rect 13920 43894 13929 43950
rect 14966 43944 15026 43946
rect 14414 43922 14474 43924
rect 13310 43775 13370 43878
rect 13862 43775 13922 43894
rect 14407 43866 14416 43922
rect 14472 43866 14481 43922
rect 14959 43888 14968 43944
rect 15024 43888 15033 43944
rect 16063 43920 16072 43976
rect 16128 43920 16137 43976
rect 17174 43970 17234 43972
rect 14414 43775 14474 43866
rect 14966 43775 15026 43888
rect 15518 43886 15578 43888
rect 15511 43830 15520 43886
rect 15576 43830 15585 43886
rect 15518 43775 15578 43830
rect 16070 43775 16130 43920
rect 17167 43914 17176 43970
rect 17232 43914 17241 43970
rect 18823 43968 18832 44024
rect 18888 43968 18897 44024
rect 17726 43938 17786 43940
rect 16622 43826 16682 43828
rect 16615 43775 16624 43826
rect 1537 43706 1546 43775
rect 1615 43770 16624 43775
rect 16680 43775 16689 43826
rect 17174 43775 17234 43914
rect 17719 43882 17728 43938
rect 17784 43882 17793 43938
rect 18278 43934 18338 43936
rect 17726 43775 17786 43882
rect 18271 43878 18280 43934
rect 18336 43878 18345 43934
rect 18278 43775 18338 43878
rect 18830 43775 18890 43968
rect 27668 43912 27728 43921
rect 27664 43854 27668 43910
rect 27728 43854 27732 43910
rect 27668 43843 27728 43852
rect 26029 43775 26098 43781
rect 28214 43775 28274 44350
rect 28766 44128 28826 44130
rect 28759 44072 28768 44128
rect 28824 44072 28833 44128
rect 28766 43775 28826 44072
rect 16680 43770 19124 43775
rect 1615 43706 19124 43770
rect 19193 43706 19204 43775
rect 26098 43706 28852 43775
rect 26029 43700 26098 43706
rect 28766 43702 28826 43706
rect 27107 43574 27173 43579
rect 27103 43518 27112 43574
rect 27168 43518 27177 43574
rect 12799 41739 12865 41745
rect 23393 41739 23459 41745
rect 27107 41739 27173 43518
rect 27670 42902 27726 42908
rect 6031 41673 12799 41739
rect 19221 41673 19227 41739
rect 19293 41673 23393 41739
rect 27101 41673 27107 41739
rect 27173 41673 27179 41739
rect 6031 41533 6097 41673
rect 12799 41667 12865 41673
rect 23393 41667 23459 41673
rect 6032 40702 6088 41533
rect 19426 40916 19482 40922
rect 27670 40916 27726 42846
rect 11000 40900 11056 40906
rect 14366 40900 19426 40916
rect 11056 40860 19426 40900
rect 23612 40860 23618 40916
rect 23674 40860 27726 40916
rect 11056 40844 14726 40860
rect 19426 40854 19482 40860
rect 11000 40838 11056 40844
rect 6032 40620 6088 40646
rect 11000 38954 11056 38992
rect 6026 38792 6032 38848
rect 6088 38792 6094 38848
rect 6032 35722 6088 38792
rect 11000 35584 11056 38898
rect 16840 6699 17040 12314
rect 19426 9824 19626 12264
rect 26162 9824 26362 9833
rect 19426 9624 26670 9824
rect 26162 9615 26362 9624
rect 16802 6690 17040 6699
rect 16802 6510 22814 6690
rect 16802 6501 16982 6510
rect 22634 4842 22814 6510
rect 26470 5450 26670 9624
rect 29570 8112 29770 12502
rect 30296 8112 30498 8118
rect 29570 7912 30498 8112
rect 30296 7903 30498 7912
rect 30296 7135 30496 7903
rect 30292 6945 30301 7135
rect 30491 6945 30500 7135
rect 30296 6940 30496 6945
rect 26470 5241 26670 5250
rect 22634 4579 22814 4662
rect -26 26 26 32
rect -26 -32 26 -26
<< via2 >>
rect 28216 44350 28272 44406
rect 7240 44108 7296 44164
rect 6688 44026 6744 44082
rect 6135 43923 6194 43982
rect 7792 43986 7848 44042
rect 8344 43906 8400 43962
rect 8896 43916 8952 43972
rect 9448 43884 9504 43940
rect 10000 43900 10056 43956
rect 10552 43874 10608 43930
rect 11104 43848 11160 43904
rect 11656 43900 11712 43956
rect 12208 43902 12264 43958
rect 12760 43910 12816 43966
rect 13312 43878 13368 43934
rect 13864 43894 13920 43950
rect 14416 43866 14472 43922
rect 14968 43888 15024 43944
rect 16072 43920 16128 43976
rect 15520 43830 15576 43886
rect 17176 43914 17232 43970
rect 18832 43968 18888 44024
rect 1546 43706 1615 43775
rect 16624 43770 16680 43826
rect 17728 43882 17784 43938
rect 18280 43878 18336 43934
rect 27668 43910 27728 43912
rect 27668 43854 27670 43910
rect 27670 43854 27726 43910
rect 27726 43854 27728 43910
rect 27668 43852 27728 43854
rect 28768 44072 28824 44128
rect 27112 43518 27168 43574
rect 30301 6945 30491 7135
rect 26470 5250 26670 5450
rect 22634 4662 22814 4842
<< metal3 >>
rect 28206 44756 28212 44820
rect 28276 44756 28282 44820
rect 27107 44614 27173 44615
rect 27102 44550 27108 44614
rect 27172 44550 27178 44614
rect 6678 44434 6684 44498
rect 6748 44434 6754 44498
rect 7230 44434 7236 44498
rect 7300 44434 7306 44498
rect 6130 44228 6199 44229
rect 6125 44161 6131 44228
rect 6198 44161 6204 44228
rect 6130 43982 6199 44161
rect 6686 44087 6746 44434
rect 7238 44169 7298 44434
rect 7235 44164 7301 44169
rect 7235 44108 7240 44164
rect 7296 44108 7301 44164
rect 7782 44150 7788 44214
rect 7852 44150 7858 44214
rect 8334 44168 8340 44232
rect 8404 44168 8410 44232
rect 8886 44174 8892 44238
rect 8956 44174 8962 44238
rect 9438 44194 9444 44258
rect 9508 44194 9514 44258
rect 9990 44220 9996 44284
rect 10060 44220 10066 44284
rect 7235 44103 7301 44108
rect 6683 44082 6749 44087
rect 6683 44026 6688 44082
rect 6744 44026 6749 44082
rect 7790 44047 7850 44150
rect 6683 44021 6749 44026
rect 7787 44042 7853 44047
rect 6130 43923 6135 43982
rect 6194 43923 6199 43982
rect 7787 43986 7792 44042
rect 7848 43986 7853 44042
rect 7787 43981 7853 43986
rect 8342 43967 8402 44168
rect 8894 43977 8954 44174
rect 8891 43972 8957 43977
rect 6130 43918 6199 43923
rect 8339 43962 8405 43967
rect 8339 43906 8344 43962
rect 8400 43906 8405 43962
rect 8891 43916 8896 43972
rect 8952 43916 8957 43972
rect 9446 43945 9506 44194
rect 9998 43961 10058 44220
rect 10542 44200 10548 44264
rect 10612 44200 10618 44264
rect 11094 44248 11100 44312
rect 11164 44248 11170 44312
rect 9995 43956 10061 43961
rect 8891 43911 8957 43916
rect 9443 43940 9509 43945
rect 8339 43901 8405 43906
rect 8342 43882 8402 43901
rect 9443 43884 9448 43940
rect 9504 43884 9509 43940
rect 9995 43900 10000 43956
rect 10056 43900 10061 43956
rect 10550 43935 10610 44200
rect 9995 43895 10061 43900
rect 10547 43930 10613 43935
rect 9443 43879 9509 43884
rect 10547 43874 10552 43930
rect 10608 43874 10613 43930
rect 11102 43909 11162 44248
rect 11646 44194 11652 44258
rect 11716 44194 11722 44258
rect 11654 43961 11714 44194
rect 12198 44176 12204 44240
rect 12268 44176 12274 44240
rect 12206 43963 12266 44176
rect 12750 44166 12756 44230
rect 12820 44166 12826 44230
rect 13302 44198 13308 44262
rect 13372 44198 13378 44262
rect 12758 43971 12818 44166
rect 12755 43966 12821 43971
rect 11651 43956 11717 43961
rect 10547 43869 10613 43874
rect 11099 43904 11165 43909
rect 11099 43848 11104 43904
rect 11160 43848 11165 43904
rect 11651 43900 11656 43956
rect 11712 43900 11717 43956
rect 11651 43895 11717 43900
rect 12203 43958 12269 43963
rect 12203 43902 12208 43958
rect 12264 43902 12269 43958
rect 12755 43910 12760 43966
rect 12816 43910 12821 43966
rect 13310 43939 13370 44198
rect 13854 44182 13860 44246
rect 13924 44182 13930 44246
rect 14406 44220 14412 44284
rect 14476 44220 14482 44284
rect 14958 44256 14964 44320
rect 15028 44256 15034 44320
rect 16062 44300 16068 44364
rect 16132 44300 16138 44364
rect 13862 43955 13922 44182
rect 13859 43950 13925 43955
rect 12755 43905 12821 43910
rect 13307 43934 13373 43939
rect 12203 43897 12269 43902
rect 13307 43878 13312 43934
rect 13368 43878 13373 43934
rect 13859 43894 13864 43950
rect 13920 43894 13925 43950
rect 14414 43927 14474 44220
rect 14966 43949 15026 44256
rect 15510 44204 15516 44268
rect 15580 44204 15586 44268
rect 14963 43944 15029 43949
rect 13859 43889 13925 43894
rect 14411 43922 14477 43927
rect 13307 43873 13373 43878
rect 14411 43866 14416 43922
rect 14472 43866 14477 43922
rect 14963 43888 14968 43944
rect 15024 43888 15029 43944
rect 15518 43891 15578 44204
rect 16070 43981 16130 44300
rect 16614 44224 16620 44288
rect 16684 44224 16690 44288
rect 16067 43976 16133 43981
rect 16067 43920 16072 43976
rect 16128 43920 16133 43976
rect 16067 43915 16133 43920
rect 14963 43883 15029 43888
rect 15515 43886 15581 43891
rect 14411 43861 14477 43866
rect 11099 43843 11165 43848
rect 11102 43824 11162 43843
rect 15515 43830 15520 43886
rect 15576 43830 15581 43886
rect 16622 43831 16682 44224
rect 17166 44198 17172 44262
rect 17236 44198 17242 44262
rect 17718 44224 17724 44288
rect 17788 44224 17794 44288
rect 17174 43975 17234 44198
rect 17171 43970 17237 43975
rect 17171 43914 17176 43970
rect 17232 43914 17237 43970
rect 17726 43943 17786 44224
rect 18270 44176 18276 44240
rect 18340 44176 18346 44240
rect 17171 43909 17237 43914
rect 17723 43938 17789 43943
rect 18278 43939 18338 44176
rect 18822 44166 18828 44230
rect 18892 44166 18898 44230
rect 18830 44029 18890 44166
rect 18827 44024 18893 44029
rect 18827 43968 18832 44024
rect 18888 43968 18893 44024
rect 18827 43963 18893 43968
rect 17723 43882 17728 43938
rect 17784 43882 17789 43938
rect 17723 43877 17789 43882
rect 18275 43934 18341 43939
rect 18275 43878 18280 43934
rect 18336 43878 18341 43934
rect 18275 43873 18341 43878
rect 15515 43825 15581 43830
rect 16619 43826 16685 43831
rect 1541 43775 1620 43780
rect 1310 43706 1316 43775
rect 1385 43706 1546 43775
rect 1615 43706 1620 43775
rect 16619 43770 16624 43826
rect 16680 43770 16685 43826
rect 16619 43765 16685 43770
rect 1541 43701 1620 43706
rect 27107 43574 27173 44550
rect 28214 44411 28274 44756
rect 28758 44744 28764 44808
rect 28828 44744 28834 44808
rect 28211 44406 28277 44411
rect 28211 44350 28216 44406
rect 28272 44350 28277 44406
rect 28211 44345 28277 44350
rect 27666 44228 27730 44240
rect 27666 44158 27730 44164
rect 27668 43917 27728 44158
rect 28766 44133 28826 44744
rect 28763 44128 28829 44133
rect 28763 44072 28768 44128
rect 28824 44072 28829 44128
rect 28763 44067 28829 44072
rect 27663 43912 27733 43917
rect 27663 43852 27668 43912
rect 27728 43852 27733 43912
rect 27663 43847 27733 43852
rect 27107 43518 27112 43574
rect 27168 43518 27173 43574
rect 27107 43513 27173 43518
rect 2709 16246 3107 16251
rect 2186 16245 3108 16246
rect 2186 16196 2709 16245
rect 254 15896 260 16196
rect 560 15896 2709 16196
rect 2186 15847 2709 15896
rect 3107 15847 3108 16245
rect 2186 15846 3108 15847
rect 2709 15841 3107 15846
rect 30296 7135 30496 7140
rect 30296 6945 30301 7135
rect 30491 6945 30496 7135
rect 30296 5955 30496 6945
rect 30291 5757 30297 5955
rect 30495 5757 30501 5955
rect 30296 5756 30496 5757
rect 26465 5450 26675 5455
rect 26465 5250 26470 5450
rect 26670 5250 26675 5450
rect 26465 5245 26675 5250
rect 22629 4842 22819 4847
rect 22629 4662 22634 4842
rect 22814 4662 22819 4842
rect 22629 4657 22819 4662
rect 22634 2546 22814 4657
rect 26470 3720 26670 5245
rect 26470 3514 26670 3520
rect 22634 2360 22814 2366
<< via3 >>
rect 28212 44756 28276 44820
rect 27108 44550 27172 44614
rect 6684 44434 6748 44498
rect 7236 44434 7300 44498
rect 6131 44161 6198 44228
rect 7788 44150 7852 44214
rect 8340 44168 8404 44232
rect 8892 44174 8956 44238
rect 9444 44194 9508 44258
rect 9996 44220 10060 44284
rect 10548 44200 10612 44264
rect 11100 44248 11164 44312
rect 11652 44194 11716 44258
rect 12204 44176 12268 44240
rect 12756 44166 12820 44230
rect 13308 44198 13372 44262
rect 13860 44182 13924 44246
rect 14412 44220 14476 44284
rect 14964 44256 15028 44320
rect 16068 44300 16132 44364
rect 15516 44204 15580 44268
rect 16620 44224 16684 44288
rect 17172 44198 17236 44262
rect 17724 44224 17788 44288
rect 18276 44176 18340 44240
rect 18828 44166 18892 44230
rect 1316 43706 1385 43775
rect 28764 44744 28828 44808
rect 27666 44164 27730 44228
rect 260 15896 560 16196
rect 2709 15847 3107 16245
rect 30297 5757 30495 5955
rect 26470 3520 26670 3720
rect 22634 2366 22814 2546
<< metal4 >>
rect 6134 44229 6194 45152
rect 6686 44499 6746 45152
rect 7238 44499 7298 45152
rect 6683 44498 6749 44499
rect 6683 44434 6684 44498
rect 6748 44434 6749 44498
rect 6683 44433 6749 44434
rect 7235 44498 7301 44499
rect 7235 44434 7236 44498
rect 7300 44434 7301 44498
rect 7235 44433 7301 44434
rect 6130 44228 6199 44229
rect 6130 44161 6131 44228
rect 6198 44161 6199 44228
rect 7790 44215 7850 45152
rect 8342 44233 8402 45152
rect 8894 44239 8954 45152
rect 9446 44259 9506 45152
rect 9998 44285 10058 45152
rect 9995 44284 10061 44285
rect 9443 44258 9509 44259
rect 8891 44238 8957 44239
rect 8339 44232 8405 44233
rect 6130 44160 6199 44161
rect 7787 44214 7853 44215
rect 6134 44152 6194 44160
rect 200 16196 600 44152
rect 7787 44150 7788 44214
rect 7852 44150 7853 44214
rect 8339 44168 8340 44232
rect 8404 44168 8405 44232
rect 8891 44174 8892 44238
rect 8956 44174 8957 44238
rect 9443 44194 9444 44258
rect 9508 44194 9509 44258
rect 9995 44220 9996 44284
rect 10060 44220 10061 44284
rect 10550 44265 10610 45152
rect 11102 44313 11162 45152
rect 11099 44312 11165 44313
rect 9995 44219 10061 44220
rect 10547 44264 10613 44265
rect 9443 44193 9509 44194
rect 8891 44173 8957 44174
rect 8339 44167 8405 44168
rect 8342 44152 8402 44167
rect 8894 44152 8954 44173
rect 9446 44152 9506 44193
rect 9998 44152 10058 44219
rect 10547 44200 10548 44264
rect 10612 44200 10613 44264
rect 11099 44248 11100 44312
rect 11164 44248 11165 44312
rect 11654 44259 11714 45152
rect 11099 44247 11165 44248
rect 11651 44258 11717 44259
rect 10547 44199 10613 44200
rect 10550 44152 10610 44199
rect 11102 44152 11162 44247
rect 11651 44194 11652 44258
rect 11716 44194 11717 44258
rect 12206 44241 12266 45152
rect 11651 44193 11717 44194
rect 12203 44240 12269 44241
rect 11654 44152 11714 44193
rect 12203 44176 12204 44240
rect 12268 44176 12269 44240
rect 12758 44231 12818 45152
rect 13310 44263 13370 45152
rect 13307 44262 13373 44263
rect 12203 44175 12269 44176
rect 12755 44230 12821 44231
rect 12206 44152 12266 44175
rect 12755 44166 12756 44230
rect 12820 44166 12821 44230
rect 13307 44198 13308 44262
rect 13372 44198 13373 44262
rect 13862 44247 13922 45152
rect 14414 44285 14474 45152
rect 14966 44321 15026 45152
rect 14963 44320 15029 44321
rect 14411 44284 14477 44285
rect 13307 44197 13373 44198
rect 13859 44246 13925 44247
rect 12755 44165 12821 44166
rect 12758 44152 12818 44165
rect 13310 44152 13370 44197
rect 13859 44182 13860 44246
rect 13924 44182 13925 44246
rect 14411 44220 14412 44284
rect 14476 44220 14477 44284
rect 14963 44256 14964 44320
rect 15028 44256 15029 44320
rect 15518 44269 15578 45152
rect 16070 44365 16130 45152
rect 16067 44364 16133 44365
rect 16067 44300 16068 44364
rect 16132 44300 16133 44364
rect 16067 44299 16133 44300
rect 14963 44255 15029 44256
rect 15515 44268 15581 44269
rect 14411 44219 14477 44220
rect 13859 44181 13925 44182
rect 13862 44152 13922 44181
rect 14414 44152 14474 44219
rect 14966 44152 15026 44255
rect 15515 44204 15516 44268
rect 15580 44204 15581 44268
rect 15515 44203 15581 44204
rect 15518 44152 15578 44203
rect 16070 44152 16130 44299
rect 16622 44289 16682 45152
rect 16619 44288 16685 44289
rect 16619 44224 16620 44288
rect 16684 44224 16685 44288
rect 17174 44263 17234 45152
rect 17726 44289 17786 45152
rect 17723 44288 17789 44289
rect 16619 44223 16685 44224
rect 17171 44262 17237 44263
rect 16622 44152 16682 44223
rect 17171 44198 17172 44262
rect 17236 44198 17237 44262
rect 17723 44224 17724 44288
rect 17788 44224 17789 44288
rect 18278 44241 18338 45152
rect 17723 44223 17789 44224
rect 18275 44240 18341 44241
rect 17171 44197 17237 44198
rect 17174 44152 17234 44197
rect 17726 44152 17786 44223
rect 18275 44176 18276 44240
rect 18340 44176 18341 44240
rect 18830 44231 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44615 27170 45152
rect 27107 44614 27173 44615
rect 27107 44550 27108 44614
rect 27172 44550 27173 44614
rect 27107 44549 27173 44550
rect 27662 44458 27722 45152
rect 28214 44821 28274 45152
rect 28211 44820 28277 44821
rect 28211 44756 28212 44820
rect 28276 44756 28277 44820
rect 28766 44809 28826 45152
rect 29318 44952 29378 45152
rect 28211 44755 28277 44756
rect 28763 44808 28829 44809
rect 28214 44746 28274 44755
rect 28763 44744 28764 44808
rect 28828 44744 28829 44808
rect 28763 44743 28829 44744
rect 27662 44372 27730 44458
rect 18275 44175 18341 44176
rect 18827 44230 18893 44231
rect 18278 44152 18338 44175
rect 18827 44166 18828 44230
rect 18892 44166 18893 44230
rect 27666 44229 27730 44372
rect 18827 44165 18893 44166
rect 27665 44228 27731 44229
rect 18830 44152 18890 44165
rect 27665 44164 27666 44228
rect 27730 44164 27731 44228
rect 27665 44163 27731 44164
rect 7787 44149 7853 44150
rect 200 15896 260 16196
rect 560 15896 600 16196
rect 200 1000 600 15896
rect 800 43775 1200 44146
rect 1315 43775 1386 43776
rect 800 43706 1316 43775
rect 1385 43706 1386 43775
rect 800 33304 1200 43706
rect 1315 43705 1386 43706
rect 800 33004 4786 33304
rect 800 1000 1200 33004
rect 2708 16245 4982 16246
rect 2708 15847 2709 16245
rect 3107 15847 4982 16245
rect 2708 15846 4982 15847
rect 30296 5955 30496 5956
rect 30296 5757 30297 5955
rect 30495 5757 30496 5955
rect 26469 3720 26671 3721
rect 26469 3520 26470 3720
rect 26670 3520 26671 3720
rect 26469 3519 26671 3520
rect 22633 2546 22815 2547
rect 22633 2366 22634 2546
rect 22814 2366 22815 2546
rect 26470 2525 26670 3519
rect 30296 2547 30496 5757
rect 22633 2333 22815 2366
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 2333
rect 26449 2323 26670 2525
rect 30295 2345 30497 2547
rect 26450 1658 26670 2323
rect 26450 936 26650 1658
rect 26450 824 26678 936
rect 26498 0 26678 824
rect 30296 656 30496 2345
rect 30296 546 30542 656
rect 30362 0 30542 546
use Mux_instance  Mux_instance_0 ~/Progetto_PISEI/mag
timestamp 1750417113
transform 1 0 3248 0 1 86
box 1148 11952 26522 35692
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel space 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 800 1000 1200 44146 0 FreeSans 1600 0 0 0 VGND
port 54 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
