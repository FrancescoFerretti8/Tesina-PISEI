magic
tech sky130A
magscale 1 2
timestamp 1749914659
<< error_p >>
rect -331 175 -269 181
rect -203 175 -141 181
rect -75 175 -13 181
rect 53 175 115 181
rect 181 175 243 181
rect 309 175 371 181
rect -331 141 -319 175
rect -203 141 -191 175
rect -75 141 -63 175
rect 53 141 65 175
rect 181 141 193 175
rect 309 141 321 175
rect -331 135 -269 141
rect -203 135 -141 141
rect -75 135 -13 141
rect 53 135 115 141
rect 181 135 243 141
rect 309 135 371 141
rect -331 -153 -269 -147
rect -203 -153 -141 -147
rect -75 -153 -13 -147
rect 53 -153 115 -147
rect 181 -153 243 -147
rect 309 -153 371 -147
rect -331 -187 -319 -153
rect -203 -187 -191 -153
rect -75 -187 -63 -153
rect 53 -187 65 -153
rect 181 -187 193 -153
rect 309 -187 321 -153
rect -331 -193 -269 -187
rect -203 -193 -141 -187
rect -75 -193 -13 -187
rect 53 -193 115 -187
rect 181 -193 243 -187
rect 309 -193 371 -187
<< nwell >>
rect -531 -325 571 313
<< pmoslvt >>
rect -335 -106 -265 94
rect -207 -106 -137 94
rect -79 -106 -9 94
rect 49 -106 119 94
rect 177 -106 247 94
rect 305 -106 375 94
<< pdiff >>
rect -393 82 -335 94
rect -393 -94 -381 82
rect -347 -94 -335 82
rect -393 -106 -335 -94
rect -265 82 -207 94
rect -265 -94 -253 82
rect -219 -94 -207 82
rect -265 -106 -207 -94
rect -137 82 -79 94
rect -137 -94 -125 82
rect -91 -94 -79 82
rect -137 -106 -79 -94
rect -9 82 49 94
rect -9 -94 3 82
rect 37 -94 49 82
rect -9 -106 49 -94
rect 119 82 177 94
rect 119 -94 131 82
rect 165 -94 177 82
rect 119 -106 177 -94
rect 247 82 305 94
rect 247 -94 259 82
rect 293 -94 305 82
rect 247 -106 305 -94
rect 375 82 433 94
rect 375 -94 387 82
rect 421 -94 433 82
rect 375 -106 433 -94
<< pdiffc >>
rect -381 -94 -347 82
rect -253 -94 -219 82
rect -125 -94 -91 82
rect 3 -94 37 82
rect 131 -94 165 82
rect 259 -94 293 82
rect 387 -94 421 82
<< nsubdiff >>
rect -495 243 -399 277
rect 439 243 535 277
rect -495 181 -461 243
rect 501 181 535 243
rect -495 -255 -461 -193
rect 501 -255 535 -193
rect -495 -289 -399 -255
rect 439 -289 535 -255
<< nsubdiffcont >>
rect -399 243 439 277
rect -495 -193 -461 181
rect 501 -193 535 181
rect -399 -289 439 -255
<< poly >>
rect -335 175 -265 191
rect -335 141 -319 175
rect -281 141 -265 175
rect -335 94 -265 141
rect -207 175 -137 191
rect -207 141 -191 175
rect -153 141 -137 175
rect -207 94 -137 141
rect -79 175 -9 191
rect -79 141 -63 175
rect -25 141 -9 175
rect -79 94 -9 141
rect 49 175 119 191
rect 49 141 65 175
rect 103 141 119 175
rect 49 94 119 141
rect 177 175 247 191
rect 177 141 193 175
rect 231 141 247 175
rect 177 94 247 141
rect 305 175 375 191
rect 305 141 321 175
rect 359 141 375 175
rect 305 94 375 141
rect -335 -153 -265 -106
rect -335 -187 -319 -153
rect -281 -187 -265 -153
rect -335 -203 -265 -187
rect -207 -153 -137 -106
rect -207 -187 -191 -153
rect -153 -187 -137 -153
rect -207 -203 -137 -187
rect -79 -153 -9 -106
rect -79 -187 -63 -153
rect -25 -187 -9 -153
rect -79 -203 -9 -187
rect 49 -153 119 -106
rect 49 -187 65 -153
rect 103 -187 119 -153
rect 49 -203 119 -187
rect 177 -153 247 -106
rect 177 -187 193 -153
rect 231 -187 247 -153
rect 177 -203 247 -187
rect 305 -153 375 -106
rect 305 -187 321 -153
rect 359 -187 375 -153
rect 305 -203 375 -187
<< polycont >>
rect -319 141 -281 175
rect -191 141 -153 175
rect -63 141 -25 175
rect 65 141 103 175
rect 193 141 231 175
rect 321 141 359 175
rect -319 -187 -281 -153
rect -191 -187 -153 -153
rect -63 -187 -25 -153
rect 65 -187 103 -153
rect 193 -187 231 -153
rect 321 -187 359 -153
<< locali >>
rect -495 243 -399 277
rect 439 243 535 277
rect -495 181 -461 243
rect 501 181 535 243
rect -335 141 -319 175
rect -281 141 -265 175
rect -207 141 -191 175
rect -153 141 -137 175
rect -79 141 -63 175
rect -25 141 -9 175
rect 49 141 65 175
rect 103 141 119 175
rect 177 141 193 175
rect 231 141 247 175
rect 305 141 321 175
rect 359 141 375 175
rect -381 82 -347 98
rect -381 -110 -347 -94
rect -253 82 -219 98
rect -253 -110 -219 -94
rect -125 82 -91 98
rect -125 -110 -91 -94
rect 3 82 37 98
rect 3 -110 37 -94
rect 131 82 165 98
rect 131 -110 165 -94
rect 259 82 293 98
rect 259 -110 293 -94
rect 387 82 421 98
rect 387 -110 421 -94
rect -335 -187 -319 -153
rect -281 -187 -265 -153
rect -207 -187 -191 -153
rect -153 -187 -137 -153
rect -79 -187 -63 -153
rect -25 -187 -9 -153
rect 49 -187 65 -153
rect 103 -187 119 -153
rect 177 -187 193 -153
rect 231 -187 247 -153
rect 305 -187 321 -153
rect 359 -187 375 -153
rect -495 -255 -461 -193
rect 501 -255 535 -193
rect -495 -289 -399 -255
rect 439 -289 535 -255
<< viali >>
rect -319 141 -281 175
rect -191 141 -153 175
rect -63 141 -25 175
rect 65 141 103 175
rect 193 141 231 175
rect 321 141 359 175
rect -381 -94 -347 82
rect -253 -94 -219 82
rect -125 -94 -91 82
rect 3 -94 37 82
rect 131 -94 165 82
rect 259 -94 293 82
rect 387 -94 421 82
rect -319 -187 -281 -153
rect -191 -187 -153 -153
rect -63 -187 -25 -153
rect 65 -187 103 -153
rect 193 -187 231 -153
rect 321 -187 359 -153
<< metal1 >>
rect -331 175 -269 181
rect -331 141 -319 175
rect -281 141 -269 175
rect -331 135 -269 141
rect -203 175 -141 181
rect -203 141 -191 175
rect -153 141 -141 175
rect -203 135 -141 141
rect -75 175 -13 181
rect -75 141 -63 175
rect -25 141 -13 175
rect -75 135 -13 141
rect 53 175 115 181
rect 53 141 65 175
rect 103 141 115 175
rect 53 135 115 141
rect 181 175 243 181
rect 181 141 193 175
rect 231 141 243 175
rect 181 135 243 141
rect 309 175 371 181
rect 309 141 321 175
rect 359 141 371 175
rect 309 135 371 141
rect -387 82 -341 94
rect -387 -94 -381 82
rect -347 -94 -341 82
rect -387 -106 -341 -94
rect -259 82 -213 94
rect -259 -94 -253 82
rect -219 -94 -213 82
rect -259 -106 -213 -94
rect -131 82 -85 94
rect -131 -94 -125 82
rect -91 -94 -85 82
rect -131 -106 -85 -94
rect -3 82 43 94
rect -3 -94 3 82
rect 37 -94 43 82
rect -3 -106 43 -94
rect 125 82 171 94
rect 125 -94 131 82
rect 165 -94 171 82
rect 125 -106 171 -94
rect 253 82 299 94
rect 253 -94 259 82
rect 293 -94 299 82
rect 253 -106 299 -94
rect 381 82 427 94
rect 381 -94 387 82
rect 421 -94 427 82
rect 381 -106 427 -94
rect -331 -153 -269 -147
rect -331 -187 -319 -153
rect -281 -187 -269 -153
rect -331 -193 -269 -187
rect -203 -153 -141 -147
rect -203 -187 -191 -153
rect -153 -187 -141 -153
rect -203 -193 -141 -187
rect -75 -153 -13 -147
rect -75 -187 -63 -153
rect -25 -187 -13 -153
rect -75 -193 -13 -187
rect 53 -153 115 -147
rect 53 -187 65 -153
rect 103 -187 115 -153
rect 53 -193 115 -187
rect 181 -153 243 -147
rect 181 -187 193 -153
rect 231 -187 243 -153
rect 181 -193 243 -187
rect 309 -153 371 -147
rect 309 -187 321 -153
rect 359 -187 371 -153
rect 309 -193 371 -187
<< properties >>
string FIXED_BBOX -478 -272 518 260
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
