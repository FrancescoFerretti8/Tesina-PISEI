** sch_path: /home/ttuser/Progetto_PISEI/xschem/parametrico.sch
**.subckt parametrico
V4 VDD GND 1.8
V5 VSS GND 0
x8 VDD VSS VSS input_only_pass output_only_pass VDD pass_gate
Vin in_only_pass VSS 1.8
Vr1 in_only_pass input_only_pass 0
.save i(vr1)
Vr2 output_only_pass net1 0
.save i(vr2)
V1 in_only_pass net1 0.01
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.option reltol=1e-5
+  abstol=1e-14
.control
  save all
  dc Vin 0.3 1.8 0.01
  let Rval = (v(input_only_pass)-v(output_only_pass))/i(Vr1)
  plot Rval
  print Rval
  op
  remzerovec
  write parametrico.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  pass_gate.sym # of pins=6
** sym_path: /home/ttuser/Progetto_PISEI/xschem/pass_gate.sym
** sch_path: /home/ttuser/Progetto_PISEI/xschem/pass_gate.sch
.subckt pass_gate VDD VSS pin Ain uscita nin
*.ipin Ain
*.ipin pin
*.ipin nin
*.ipin VDD
*.ipin VSS
*.opin uscita
XM2 Ain nin uscita VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 uscita pin Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=16 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
