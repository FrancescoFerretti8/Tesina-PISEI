magic
tech sky130A
magscale 1 2
timestamp 1749982881
<< error_p >>
rect -269 172 -211 178
rect -77 172 -19 178
rect 115 172 173 178
rect 307 172 365 178
rect -269 138 -257 172
rect -77 138 -65 172
rect 115 138 127 172
rect 307 138 319 172
rect -269 132 -211 138
rect -77 132 -19 138
rect 115 132 173 138
rect 307 132 365 138
rect -365 -138 -307 -132
rect -173 -138 -115 -132
rect 19 -138 77 -132
rect 211 -138 269 -132
rect -365 -172 -353 -138
rect -173 -172 -161 -138
rect 19 -172 31 -138
rect 211 -172 223 -138
rect -365 -178 -307 -172
rect -173 -178 -115 -172
rect 19 -178 77 -172
rect 211 -178 269 -172
<< pwell >>
rect -551 -310 551 310
<< nmoslvt >>
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
<< ndiff >>
rect -413 88 -351 100
rect -413 -88 -401 88
rect -367 -88 -351 88
rect -413 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 413 100
rect 351 -88 367 88
rect 401 -88 413 88
rect 351 -100 413 -88
<< ndiffc >>
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
<< psubdiff >>
rect -515 240 -419 274
rect 419 240 515 274
rect -515 178 -481 240
rect 481 178 515 240
rect -515 -240 -481 -178
rect 481 -240 515 -178
rect -515 -274 -419 -240
rect 419 -274 515 -240
<< psubdiffcont >>
rect -419 240 419 274
rect -515 -178 -481 178
rect 481 -178 515 178
rect -419 -274 419 -240
<< poly >>
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 321 100 351 122
rect -351 -122 -321 -100
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
<< polycont >>
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
<< locali >>
rect -515 240 -419 274
rect 419 240 515 274
rect -515 178 -481 240
rect 481 178 515 240
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect -515 -240 -481 -178
rect 481 -240 515 -178
rect -515 -274 -419 -240
rect 419 -274 515 -240
<< viali >>
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
<< metal1 >>
rect -269 172 -211 178
rect -269 138 -257 172
rect -223 138 -211 172
rect -269 132 -211 138
rect -77 172 -19 178
rect -77 138 -65 172
rect -31 138 -19 172
rect -77 132 -19 138
rect 115 172 173 178
rect 115 138 127 172
rect 161 138 173 172
rect 115 132 173 138
rect 307 172 365 178
rect 307 138 319 172
rect 353 138 365 172
rect 307 132 365 138
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect -365 -138 -307 -132
rect -365 -172 -353 -138
rect -319 -172 -307 -138
rect -365 -178 -307 -172
rect -173 -138 -115 -132
rect -173 -172 -161 -138
rect -127 -172 -115 -138
rect -173 -178 -115 -172
rect 19 -138 77 -132
rect 19 -172 31 -138
rect 65 -172 77 -138
rect 19 -178 77 -172
rect 211 -138 269 -132
rect 211 -172 223 -138
rect 257 -172 269 -138
rect 211 -178 269 -172
<< properties >>
string FIXED_BBOX -498 -257 498 257
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
