** sch_path: /home/ttuser/tt10-analog-buffer/xschem/testbenchtwo.sch
**.subckt testbenchtwo OUT
*.opin OUT
x1 VDD VSS net1 in buffer_casa
V2 VDD GND 1.8
V3 VSS GND 0
V1 in GND pwl 0 0 10n 0 10.1n 1.8 20n 1.8 20.1n 0
R2 OUT net1 500 m=1
C1 net1 VSS 5p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.control
tran 100p 50n
write testbenchtwo.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  buffer_casa.sym # of pins=4
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/buffer_casa.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/buffer_casa.sch
.subckt buffer_casa VDD VSS OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 outm IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outm IN VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT outm VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT outm VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
