** sch_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sch
.subckt pass_gate Inp VDD out Ain VSS Inn
*.PININFO Inp:I Inn:I out:O Ain:I VDD:I VSS:I
XM10 out Inp Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=32 nf=32 m=1
XM1 Ain Inn out VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=16 nf=16 m=1
.ends
.end
