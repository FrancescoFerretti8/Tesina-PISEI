magic
tech sky130A
magscale 1 2
timestamp 1750417113
<< metal1 >>
rect 11754 30998 11874 31004
rect 11874 30878 13220 30998
rect 11754 30872 11874 30878
rect 13100 29374 13220 30878
rect 22920 30154 23120 30160
rect 15466 29374 16713 29379
rect 13100 29254 16713 29374
rect 15466 29225 16713 29254
rect 22920 29200 23120 29954
rect 11274 29094 11394 29100
rect 11394 28974 12578 29094
rect 11274 28968 11394 28974
rect 11392 27070 11398 27190
rect 11518 27070 11524 27190
rect 10784 25286 10904 25292
rect 10784 21062 10904 25166
rect 11398 23728 11518 27070
rect 12458 26576 12578 28974
rect 15678 28797 15878 28803
rect 15878 28597 16666 28797
rect 15678 28591 15878 28597
rect 12710 28072 12830 28078
rect 15466 28072 16519 28085
rect 12830 27952 16519 28072
rect 12710 27946 12830 27952
rect 15466 27934 16519 27952
rect 15466 26576 16543 26589
rect 12458 26456 16543 26576
rect 15466 26427 16543 26456
rect 16448 25793 16454 25993
rect 16654 25793 16660 25993
rect 15466 25276 16600 25278
rect 14058 25156 14064 25276
rect 14184 25158 16600 25276
rect 14184 25156 15518 25158
rect 24312 24311 25896 24511
rect 26096 24311 26102 24511
rect 15466 23728 16610 23750
rect 11398 23608 16610 23728
rect 15466 23602 16610 23608
rect 14758 22426 14878 22432
rect 15466 22426 16494 22434
rect 14878 22314 16494 22426
rect 14878 22306 15502 22314
rect 14758 22300 14878 22306
rect 15466 21062 16778 21087
rect 10784 20942 16778 21062
rect 15466 20914 16778 20942
rect 15466 19796 16552 19804
rect 15184 19684 16552 19796
rect 15184 19676 15474 19684
rect 15184 18420 15304 19676
rect 23424 18578 23624 19081
rect 15178 18300 15184 18420
rect 15304 18300 15310 18420
rect 23364 18084 23664 18578
rect 23358 17784 23670 18084
rect 16742 16072 16937 16078
rect 23404 16072 23599 17784
rect 16937 15877 23599 16072
rect 16742 15871 16937 15877
<< via1 >>
rect 11754 30878 11874 30998
rect 22920 29954 23120 30154
rect 11274 28974 11394 29094
rect 11398 27070 11518 27190
rect 10784 25166 10904 25286
rect 15678 28597 15878 28797
rect 12710 27952 12830 28072
rect 16454 25793 16654 25993
rect 14064 25156 14184 25276
rect 25896 24311 26096 24511
rect 14758 22306 14878 22426
rect 15184 18300 15304 18420
rect 16742 15877 16937 16072
<< metal2 >>
rect 2784 31904 2840 35692
rect 7752 31954 7808 35692
rect 14445 32986 14454 33186
rect 14654 32986 23120 33186
rect 10029 30998 10139 31002
rect 10024 30993 11754 30998
rect 10024 30883 10029 30993
rect 10139 30883 11754 30993
rect 10024 30878 11754 30883
rect 11874 30878 11880 30998
rect 10029 30874 10139 30878
rect 22920 30154 23120 32986
rect 22914 29954 22920 30154
rect 23120 29954 23126 30154
rect 9985 29094 10095 29098
rect 9980 29089 11274 29094
rect 9980 28979 9985 29089
rect 10095 28979 11274 29089
rect 9980 28974 11274 28979
rect 11394 28974 11400 29094
rect 9985 28970 10095 28974
rect 15672 28597 15678 28797
rect 15878 28597 15884 28797
rect 12704 27952 12710 28072
rect 12830 27952 12836 28072
rect 10103 27190 10213 27194
rect 11398 27190 11518 27196
rect 10098 27185 11398 27190
rect 10098 27075 10103 27185
rect 10213 27075 11398 27185
rect 10098 27070 11398 27075
rect 10103 27066 10213 27070
rect 11398 27064 11518 27070
rect 10091 25286 10201 25290
rect 10086 25281 10784 25286
rect 10086 25171 10091 25281
rect 10201 25171 10784 25281
rect 10086 25166 10784 25171
rect 10904 25166 10910 25286
rect 10091 25162 10201 25166
rect 12710 25001 12830 27952
rect 14064 25276 14184 25282
rect 12706 24891 12715 25001
rect 12825 24891 12834 25001
rect 12710 24886 12830 24891
rect 14064 22973 14184 25156
rect 14060 22863 14069 22973
rect 14179 22863 14188 22973
rect 14064 22858 14184 22863
rect 14752 22306 14758 22426
rect 14878 22306 14884 22426
rect 14758 20365 14878 22306
rect 14754 20255 14763 20365
rect 14873 20255 14882 20365
rect 14758 20250 14878 20255
rect 15184 18420 15304 18426
rect 12131 17670 12241 17674
rect 15184 17670 15304 18300
rect 12126 17665 15304 17670
rect 12126 17555 12131 17665
rect 12241 17555 15304 17665
rect 12126 17550 15304 17555
rect 12131 17546 12241 17550
rect 13592 16906 15188 16916
rect 15678 16906 15878 28597
rect 16454 25993 16654 25999
rect 13592 16716 15878 16906
rect 13592 14007 13792 16716
rect 15088 16706 15878 16716
rect 16178 25793 16454 25993
rect 13588 13817 13796 14007
rect 13592 12028 13792 13817
rect 16178 11952 16378 25793
rect 16454 25787 16654 25793
rect 25896 24511 26096 24517
rect 26096 24311 26522 24511
rect 25896 24305 26096 24311
rect 16747 16072 16932 16076
rect 16736 15877 16742 16072
rect 16937 15877 16943 16072
rect 16747 15873 16932 15877
rect 26322 12080 26522 24311
<< via2 >>
rect 14454 32986 14654 33186
rect 10029 30883 10139 30993
rect 9985 28979 10095 29089
rect 10103 27075 10213 27185
rect 10091 25171 10201 25281
rect 12715 24891 12825 25001
rect 14069 22863 14179 22973
rect 14763 20255 14873 20365
rect 12131 17555 12241 17665
rect 16747 15882 16932 16067
<< metal3 >>
rect 14449 33186 14659 33191
rect 10300 32986 10306 33186
rect 10506 32986 14454 33186
rect 14654 32986 14659 33186
rect 14449 32981 14659 32986
rect 10024 30993 10144 30998
rect 10024 30883 10029 30993
rect 10139 30883 10144 30993
rect 10024 30878 10144 30883
rect 9980 29089 10100 29094
rect 9980 28979 9985 29089
rect 10095 28979 10100 29089
rect 9980 28974 10100 28979
rect 10098 27185 10218 27190
rect 10098 27075 10103 27185
rect 10213 27075 10218 27185
rect 10098 27070 10218 27075
rect 10086 25281 10206 25286
rect 10086 25171 10091 25281
rect 10201 25171 10206 25281
rect 10086 25166 10206 25171
rect 12710 25001 12830 25006
rect 12710 24891 12715 25001
rect 12825 24891 12830 25001
rect 12710 23382 12830 24891
rect 10106 23262 12830 23382
rect 14064 22973 14184 22978
rect 14064 22863 14069 22973
rect 14179 22863 14184 22973
rect 14064 21478 14184 22863
rect 10142 21358 14184 21478
rect 14758 20365 14878 20370
rect 14758 20255 14763 20365
rect 14873 20255 14878 20365
rect 14758 19574 14878 20255
rect 10044 19454 14878 19574
rect 9998 17665 12246 17670
rect 9998 17555 12131 17665
rect 12241 17555 12246 17665
rect 9998 17550 12246 17555
rect 9513 16124 9750 16130
rect 9512 15855 9513 16094
rect 9750 16072 11217 16094
rect 9750 16067 16937 16072
rect 9750 15882 16747 16067
rect 16932 15882 16937 16067
rect 9750 15877 16937 15882
rect 9750 15855 11217 15877
rect 9513 15818 9750 15824
<< via3 >>
rect 10306 32986 10506 33186
rect 9513 15824 9750 16124
<< metal4 >>
rect 1148 33208 9682 33218
rect 10425 33208 10627 33209
rect 1148 33186 10627 33208
rect 1148 33008 10306 33186
rect 1148 32918 9682 33008
rect 10305 32986 10306 33008
rect 10506 33007 10627 33186
rect 10506 32986 10507 33007
rect 10305 32985 10507 32986
rect 3114 30942 3414 32918
rect 5086 30960 5386 32918
rect 7068 30914 7368 32918
rect 9042 30924 9342 32918
rect 2124 16124 2424 17454
rect 4098 16124 4398 17482
rect 6082 16124 6382 17482
rect 8058 16124 8358 17482
rect 9449 16124 9751 16125
rect 1184 15824 9513 16124
rect 9750 15824 9751 16124
rect 9449 15823 9751 15824
use Decoder  Decoder_0
timestamp 1750082308
transform 1 0 282 0 -1 32094
box 974 0 10000 14736
use Mux  Mux_0
timestamp 1750003929
transform 1 0 17666 0 1 28199
box -1260 -9331 6846 1730
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
