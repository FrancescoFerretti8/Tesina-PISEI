** sch_path: /home/ttuser/tt10-analog-buffer/xschem/untitled-3.sch
.subckt untitled-3

x1 net1 net3 net4 net5 net6 net7 net8 net9 net10 net11 net12 net13 Mux
.ends

* expanding   symbol:  Mux.sym # of pins=14
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/Mux.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/Mux.sch
.subckt Mux VDD VSS n0 A0 p0 n1 A1 p1 n2 p2 n3 OUT
*.PININFO OUT:O n0:I p0:I n1:I p1:I VSS:I VDD:I VDD:I A0:I A1:I n2:I n3:I p2:I p2:I
x1 n0 VDD OUT A0 VSS p0 pass_gate
x2 n1 VDD OUT A1 VSS p1 pass_gate
x3 n2 VDD OUT VDD VSS p2 pass_gate
x4 n3 VDD OUT net1 VSS p2 pass_gate
R6 net1 VDD 500 m=1
R7 GND net1 500 m=1
.ends


* expanding   symbol:  pass_gate.sym # of pins=6
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sch
.subckt pass_gate Inp VDD out Ain VSS Inn
*.PININFO Inp:I Inn:I out:O Ain:I VDD:I VSS:I
XM10 out Inp Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=32 nf=32 m=1
XM1 Ain Inn out VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=16 nf=16 m=1
.ends

.GLOBAL GND
.end
