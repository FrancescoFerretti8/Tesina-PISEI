** sch_path: /home/ttuser/Progetto_PISEI/xschem/PISEI_test.sch
**.subckt PISEI_test Uscita
*.opin Uscita
V4 VDD GND 1.8
V5 VSS GND 0
V2 net3 VSS sin(0.9 0.7 10Meg 0 0 0)
V3 net1 VSS pwl 10n 0 20n 1.8 80n 1.8 90n 0 500n 0
V1 a VSS pwl 100n 0 100.1n 1.8 200n 1.8 200.1n 0 300n 0 300.1n 1.8 400n 1.8 400.1n 0 500n 0
V6 b VSS pwl 200n 0 200.1n 1.8 400n 1.8 400.1n 0 500n 0
x2 VSS net1 input0 pad_model
x3 VSS net3 input2 pad_model
x4 VSS net2 Uscita pad_model
x1 b input2 input0 net2 a VSS VDD test_pisei_parax
**** begin user architecture code



.option reltol=1e-5
+  abstol=1e-14 savecurrents
.control
  save all
  op
  remzerovec
write PISEI_test.raw
set appendwrite
tran 100n 500n
write PISEI_test.raw
set appendwrite
*ac dec 10 1 1e12
*write PISEI_test.raw
*set appendwrite
.endc




** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  pad_model.sym # of pins=3
** sym_path: /home/ttuser/Progetto_PISEI/xschem/pad_model.sym
** sch_path: /home/ttuser/Progetto_PISEI/xschem/pad_model.sch
.subckt pad_model VGND pin mod
*.iopin pin
*.iopin mod
*.iopin VGND
C1 pin VGND 2p m=1
V1 VAPWR VGND 3.3
R1 net1 pin 1 m=1
L1 net2 net1 1n m=1
C2 net2 VGND 3p m=1
R2 net3 net2 50 m=1
C3 mod VGND 250f m=1
XM5 net3 VGND mod VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 VAPWR VGND VAPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net3 VGND VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net3 VAPWR mod VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  test_pisei_parax.sym # of pins=7
** sym_path: /home/ttuser/Progetto_PISEI/xschem/test_pisei_parax.sym
.include /home/ttuser/Progetto_PISEI/mag/test_PISEI.sim.spice
.GLOBAL GND
.end
