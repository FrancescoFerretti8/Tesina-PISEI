** sch_path: /home/ttuser/tt10-analog-buffer/xschem/Mux_per_magic.sch
.subckt Mux_per_magic

x1 net1 net2 net3 net4 net5 net6 net7 net8 net9 net10 net11 net12 net13 net14 net15 Mux
.ends

* expanding   symbol:  Mux.sym # of pins=15
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/Mux.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/Mux.sch
.subckt Mux VDD out VSS n0 A0 p0 n1 A1 p1 n2 A2 p2 n3 A3 p3
*.PININFO VDD:I VSS:I A0:I n0:I p0:I out:I A1:I n1:I p1:I A2:I n2:I p2:I A3:I n3:I p3:I
x1 n0 VDD out A0 VSS p0 pass_gate
x2 n1 VDD out A1 VSS p1 pass_gate
x3 n2 VDD out A2 VSS p2 pass_gate
x4 n3 VDD out A3 VSS p3 pass_gate
.ends


* expanding   symbol:  pass_gate.sym # of pins=6
** sym_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sym
** sch_path: /home/ttuser/tt10-analog-buffer/xschem/pass_gate.sch
.subckt pass_gate Inp VDD out Ain VSS Inn
*.PININFO Inp:I Inn:I out:O Ain:I VDD:I VSS:I
XM10 out Inp Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=32 nf=32 m=1
XM1 Ain Inn out VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=16 nf=16 m=1
.ends

.end
