* NGSPICE file created from Decoder_parax.ext - technology: sky130A

.subckt Decoder_parax VGND n[0] n[1] n[2] p[0] a p[3] p[1] p[2] n[3] b VPWR
X0 VGND.t201 VPWR.t218 VGND.t200 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1 n[0].t3 net2 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_4903_5263# net1 VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t96 VGND.t216 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4 VPWR.t42 a_2879_2223# n[1].t7 VPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5 a_2557_2767# net2 VPWR.t128 VPWR.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_4903_5263# net2 p[3].t3 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 n[3].t7 a_5179_2223# VPWR.t210 VPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 p[1].t3 a_5179_2767# VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t198 VPWR.t219 VGND.t197 VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X10 VGND.t24 a_2879_2223# n[1].t3 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 VPWR.t81 a_4075_2767# n[2].t7 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 n[3].t3 a_5179_2223# VGND.t215 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND.t196 VPWR.t220 VGND.t195 VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X14 VPWR.t126 net2 a_2557_2767# VPWR.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t193 VPWR.t221 VGND.t192 VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X16 VPWR.t98 VGND.t217 VPWR.t97 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X17 VPWR.t5 _04_ a_5179_2767# VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X18 a_4903_5263# net2 p[3].t2 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND.t190 VPWR.t222 VGND.t189 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X20 a_3523_2767# net2 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VPWR.t157 VGND.t218 VPWR.t156 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X22 VPWR.t209 a_5179_2223# n[3].t6 VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X23 VGND.t30 a_5179_2767# p[1].t2 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VGND.t112 net1 a_4819_2883# VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 p[3].t7 net2 VPWR.t124 VPWR.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t110 net1 a_4837_3339# VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 n[2].t6 a_4075_2767# VPWR.t79 VPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X28 VPWR.t159 VGND.t219 VPWR.t158 VPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X29 VGND.t213 a_5179_2223# n[3].t2 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 p[2].t7 a_5179_4399# VPWR.t19 VPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X31 VGND.t120 _05_ a_5179_4399# VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X32 p[0].t7 a_5179_3311# VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X33 n[0].t11 net1 a_2557_2767# VPWR.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 VGND.t188 VPWR.t223 VGND.t187 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X35 _04_ a_4819_2883# VGND.t42 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X36 VGND.t186 VPWR.t224 VGND.t185 VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X37 VPWR.t198 _01_ a_4075_2767# VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X38 p[0].t3 a_5179_3311# VGND.t118 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X39 VPWR.t77 a_4075_2767# n[2].t5 VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X40 VPWR.t8 VGND.t220 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X41 VGND.t77 _00_ a_2879_2223# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X42 VPWR.t17 a_5179_4399# p[2].t6 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X43 n[2].t3 a_4075_2767# VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X44 VPWR.t192 a_5179_3311# p[0].t6 VPWR.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X45 a_5095_5737# a_4903_5493# VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X46 VPWR.t11 VGND.t221 VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X47 n[0].t10 net1 a_2557_2767# VPWR.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X48 VPWR.t203 VGND.t222 VPWR.t202 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X49 VGND.t61 net2 a_4760_2473# VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VGND.t117 a_5179_3311# p[0].t2 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X51 VPWR.t184 net1 p[3].t11 VPWR.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X52 VPWR.t206 VGND.t223 VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X53 VGND.t184 VPWR.t225 VGND.t183 VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X54 a_4837_3339# net2 a_4751_3339# VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X55 VGND.t181 VPWR.t226 VGND.t180 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X56 VPWR.t214 VGND.t224 VPWR.t213 VPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X57 VGND.t108 net1 a_3793_3133# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X58 p[2].t5 a_5179_4399# VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X59 VGND.t178 VPWR.t227 VGND.t177 VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X60 VGND.t38 a_4075_2767# n[2].t2 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X61 VPWR.t154 a_2327_5487# net1 VPWR.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X62 VPWR.t217 VGND.t225 VPWR.t216 VPWR.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X63 p[0].t5 a_5179_3311# VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X64 VGND.t176 VPWR.t228 VGND.t175 VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X65 VGND.t106 net1 a_4903_5263# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X66 VPWR.t122 net2 a_2557_2767# VPWR.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X67 p[0].t1 a_5179_3311# VGND.t116 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X68 net2 a_4312_5461# VPWR.t163 VPWR.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X69 VPWR.t182 net1 p[3].t10 VPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X70 VGND.t173 VPWR.t229 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X71 VPWR.t150 _02_ a_5179_2223# VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X72 VPWR.t13 a_5179_4399# p[2].t4 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X73 VPWR.t120 net2 p[3].t6 VPWR.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X74 VPWR.t91 VGND.t226 VPWR.t90 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X75 n[2].t1 a_4075_2767# VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X76 VPWR.t93 VGND.t227 VPWR.t92 VPWR.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X77 VPWR.t188 a_5179_3311# p[0].t4 VPWR.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X78 VGND.t58 net2 a_4627_3127# VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X79 VGND.t105 net1 n[0].t7 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X80 VPWR.t56 VGND.t228 VPWR.t55 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X81 VPWR.t59 VGND.t229 VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X82 p[2].t3 a_5179_4399# VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X83 VPWR.t51 VGND.t230 VPWR.t50 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X84 VPWR.t180 net1 a_3703_2767# VPWR.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X85 VGND.t115 a_5179_3311# p[0].t0 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X86 a_3793_3133# a_3523_2767# a_3703_2767# VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X87 p[3].t1 net2 a_4903_5263# VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X88 _01_ a_3703_2767# VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X89 VGND.t170 VPWR.t230 VGND.t169 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X90 _02_ a_4751_3339# VPWR.t130 VPWR.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X91 VPWR.t118 net2 p[3].t5 VPWR.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X92 VGND.t167 VPWR.t231 VGND.t166 VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X93 VGND.t87 a_4312_5461# net2 VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X94 VGND.t34 a_4075_2767# n[2].t0 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X95 VGND.t164 VPWR.t232 VGND.t163 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X96 VGND.t44 a.t0 a_2327_5487# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X97 VPWR.t116 net2 a_2599_3677# VPWR.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X98 VGND.t103 net1 n[0].t6 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X99 VGND.t11 a_5179_4399# p[2].t2 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X100 a_4312_5461# b.t0 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X101 VPWR.t53 VGND.t231 VPWR.t52 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X102 _03_ a_4760_2473# VPWR.t132 VPWR.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X103 a_4901_2883# a_4627_3127# a_4819_2883# VPWR.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X104 net1 a_2327_5487# VGND.t83 VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X105 _05_ a_5095_5737# VGND.t73 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X106 VPWR.t100 a.t1 a_2327_5487# VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X107 VPWR.t28 VGND.t232 VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X108 a_4819_2883# a_4627_3127# VGND.t207 VGND.t206 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X109 VPWR.t30 VGND.t233 VPWR.t29 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X110 _04_ a_4819_2883# VPWR.t89 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X111 a_4312_5461# b.t1 VPWR.t212 VPWR.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X112 a_5177_5737# a_4903_5493# a_5095_5737# VPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X113 VGND.t162 VPWR.t233 VGND.t161 VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X114 p[2].t1 a_5179_4399# VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X115 VGND.t55 net2 a_5095_5737# VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X116 a_4842_2473# net1 a_4760_2473# VPWR.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X117 VPWR.t114 net2 a_3523_2767# VPWR.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X118 VGND.t53 net2 n[0].t2 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X119 VGND.t159 VPWR.t234 VGND.t158 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X120 VGND.t157 VPWR.t235 VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X121 VGND.t101 net1 a_4903_5263# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X122 VPWR.t70 VGND.t234 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X123 VGND.t3 _04_ a_5179_2767# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X124 p[1].t7 a_5179_2767# VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X125 VPWR.t196 _05_ a_5179_4399# VPWR.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X126 VGND.t154 VPWR.t236 VGND.t153 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X127 VGND.t152 VPWR.t237 VGND.t151 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X128 VPWR.t34 _03_ a_5179_3311# VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X129 VGND.t7 a_5179_4399# p[2].t0 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X130 VGND.t79 _02_ a_5179_2223# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X131 VPWR.t177 net1 a_4901_2883# VPWR.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X132 VPWR.t73 VGND.t235 VPWR.t72 VPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X133 VGND.t51 net2 n[0].t1 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X134 VGND.t149 VPWR.t238 VGND.t148 VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X135 p[3].t9 net1 VPWR.t175 VPWR.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X136 _00_ a_2599_3677# VPWR.t200 VPWR.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X137 a_4760_2473# net1 VGND.t99 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X138 VGND.t146 VPWR.t239 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X139 VPWR.t84 VGND.t236 VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X140 VPWR.t65 a_5179_2767# p[1].t6 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X141 VPWR.t87 VGND.t237 VPWR.t86 VPWR.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X142 VPWR.t173 net1 a_4751_3339# VPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X143 VGND.t49 net2 a_2689_3311# VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X144 VGND.t203 _01_ a_4075_2767# VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X145 VPWR.t112 net2 a_5177_5737# VPWR.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 VPWR.t146 VGND.t238 VPWR.t145 VPWR.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X147 VGND.t143 VPWR.t240 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X148 _02_ a_4751_3339# VGND.t69 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X149 VGND.t140 VPWR.t241 VGND.t139 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X150 n[0].t0 net2 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 a_2557_2767# net1 n[0].t9 VPWR.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X152 p[3].t0 net2 a_4903_5263# VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X153 VPWR.t149 VGND.t239 VPWR.t148 VPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X154 a_2419_3677# net1 VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X155 p[1].t5 a_5179_2767# VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X156 VPWR.t140 VGND.t240 VPWR.t139 VPWR.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X157 p[3].t4 net2 VPWR.t104 VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X158 n[1].t6 a_2879_2223# VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X159 _01_ a_3703_2767# VPWR.t32 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X160 VGND.t95 net1 a_4903_5493# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 _03_ a_4760_2473# VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X162 VGND.t137 VPWR.t242 VGND.t136 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X163 VPWR.t143 VGND.t241 VPWR.t142 VPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X164 n[0].t5 net1 VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X165 VGND.t134 VPWR.t243 VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X166 VPWR.t45 VGND.t242 VPWR.t44 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X167 n[1].t2 a_2879_2223# VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X168 VPWR.t48 VGND.t243 VPWR.t47 VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X169 a_2557_2767# net1 n[0].t8 VPWR.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_2689_3311# a_2419_3677# a_2599_3677# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X171 VPWR.t61 a_5179_2767# p[1].t4 VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X172 VGND.t81 a_2327_5487# net1 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X173 a_3703_2767# a_3523_2767# VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X174 VGND.t131 VPWR.t244 VGND.t130 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X175 a_4751_3339# net2 VPWR.t110 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X176 VPWR.t38 a_2879_2223# n[1].t5 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X177 n[3].t5 a_5179_2223# VPWR.t208 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X178 p[1].t1 a_5179_2767# VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X179 net2 a_4312_5461# VGND.t85 VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X180 VGND.t20 a_2879_2223# n[1].t1 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X181 n[0].t4 net1 VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X182 VPWR.t169 net1 a_2419_3677# VPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X183 a_2599_3677# a_2419_3677# VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X184 n[3].t1 a_5179_2223# VGND.t211 VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X185 VGND.t128 VPWR.t245 VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X186 VGND.t125 VPWR.t246 VGND.t124 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X187 a_4903_5263# net1 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 VPWR.t137 _00_ a_2879_2223# VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X189 VGND.t16 _03_ a_5179_3311# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X190 VPWR.t161 a_4312_5461# net2 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X191 a_4903_5493# net1 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X192 VPWR.t22 VGND.t244 VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X193 a_2557_2767# net2 VPWR.t108 VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X194 n[1].t4 a_2879_2223# VPWR.t36 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X195 a_4627_3127# net2 VPWR.t106 VPWR.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 p[3].t8 net1 VPWR.t165 VPWR.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 VPWR.t207 a_5179_2223# n[3].t4 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X198 VGND.t26 a_5179_2767# p[1].t0 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 VGND.t123 VPWR.t247 VGND.t122 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X200 VPWR.t25 VGND.t245 VPWR.t24 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X201 _00_ a_2599_3677# VGND.t205 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X202 n[2].t4 a_4075_2767# VPWR.t75 VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X203 net1 a_2327_5487# VPWR.t152 VPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X204 _05_ a_5095_5737# VPWR.t134 VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X205 n[1].t0 a_2879_2223# VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X206 VPWR.t102 net2 a_4842_2473# VPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X207 VGND.t209 a_5179_2223# n[3].t0 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 VPWR VPWR.t155 1719.47
R1 VPWR.t155 VPWR 1547.82
R2 VPWR VPWR.t68 975.178
R3 VPWR VPWR.t85 975.178
R4 VPWR.t68 VPWR 877.827
R5 VPWR.t85 VPWR 877.827
R6 VPWR.t26 VPWR.t71 816.822
R7 VPWR.n122 VPWR.t25 812.014
R8 VPWR.n20 VPWR.t84 804.731
R9 VPWR.n23 VPWR.t91 804.731
R10 VPWR.n497 VPWR.t87 804.731
R11 VPWR.n483 VPWR.t86 804.731
R12 VPWR.n497 VPWR.t93 804.731
R13 VPWR.n483 VPWR.t92 804.731
R14 VPWR.n442 VPWR.t70 804.731
R15 VPWR.n46 VPWR.t69 804.731
R16 VPWR.n442 VPWR.t214 804.731
R17 VPWR.n46 VPWR.t213 804.731
R18 VPWR.t10 VPWR.n39 804.731
R19 VPWR.n696 VPWR.t205 804.731
R20 VPWR.n501 VPWR.t45 804.731
R21 VPWR.n504 VPWR.t53 804.731
R22 VPWR.n571 VPWR.t51 804.731
R23 VPWR.n534 VPWR.t50 804.731
R24 VPWR.n532 VPWR.t149 804.731
R25 VPWR.n536 VPWR.t217 804.731
R26 VPWR.n141 VPWR.t148 804.731
R27 VPWR.n136 VPWR.t216 804.731
R28 VPWR.n93 VPWR.t24 804.731
R29 VPWR.n80 VPWR.t56 804.731
R30 VPWR.n83 VPWR.t98 804.731
R31 VPWR.n575 VPWR.t30 804.731
R32 VPWR.n578 VPWR.t8 804.731
R33 VPWR.n646 VPWR.t146 804.731
R34 VPWR.n160 VPWR.t145 804.731
R35 VPWR.n185 VPWR.t159 804.731
R36 VPWR.n188 VPWR.t143 804.731
R37 VPWR.n608 VPWR.t203 804.731
R38 VPWR.n611 VPWR.t22 804.731
R39 VPWR.n403 VPWR.t157 804.731
R40 VPWR.n378 VPWR.t156 804.731
R41 VPWR.t215 VPWR.t147 772.086
R42 VPWR.n41 VPWR.t10 751.692
R43 VPWR.t205 VPWR.n695 751.692
R44 VPWR.t84 VPWR.n19 725.173
R45 VPWR.t91 VPWR.n22 725.173
R46 VPWR.t45 VPWR.n500 725.173
R47 VPWR.t53 VPWR.n503 725.173
R48 VPWR.t56 VPWR.n79 725.173
R49 VPWR.t98 VPWR.n82 725.173
R50 VPWR.t30 VPWR.n574 725.173
R51 VPWR.t8 VPWR.n577 725.173
R52 VPWR.t159 VPWR.n184 725.173
R53 VPWR.t143 VPWR.n187 725.173
R54 VPWR.t203 VPWR.n607 725.173
R55 VPWR.t22 VPWR.n610 725.173
R56 VPWR.n344 VPWR.t167 701.529
R57 VPWR.n166 VPWR.t106 701.014
R58 VPWR.n115 VPWR.t110 671.408
R59 VPWR VPWR.t94 636.293
R60 VPWR.n197 VPWR.n194 604.076
R61 VPWR.n197 VPWR.n195 604.076
R62 VPWR.n636 VPWR.n268 603.106
R63 VPWR.n32 VPWR.n17 599.808
R64 VPWR.n71 VPWR.n70 599.808
R65 VPWR.n242 VPWR.n159 599.808
R66 VPWR.n591 VPWR.n570 599.159
R67 VPWR.n260 VPWR.n153 599.159
R68 VPWR.n562 VPWR.n530 585
R69 VPWR.n564 VPWR.n563 585
R70 VPWR.n251 VPWR.n250 585
R71 VPWR.n253 VPWR.n252 585
R72 VPWR.t166 VPWR.t135 568.225
R73 VPWR VPWR.t138 494.238
R74 VPWR.t162 VPWR 461.683
R75 VPWR.t94 VPWR 458.724
R76 VPWR.t57 VPWR 414.577
R77 VPWR.t46 VPWR 414.577
R78 VPWR.t12 VPWR.t82 404.505
R79 VPWR.t60 VPWR.t141 404.505
R80 VPWR.n693 VPWR.t206 389.521
R81 VPWR.n43 VPWR.t11 389.361
R82 VPWR.n666 VPWR.t59 388.656
R83 VPWR.n274 VPWR.t47 388.656
R84 VPWR.n605 VPWR.t48 388.656
R85 VPWR.n369 VPWR.t95 388.656
R86 VPWR.n372 VPWR.t96 388.656
R87 VPWR.n123 VPWR.t58 385.026
R88 VPWR.n418 VPWR.t139 381.443
R89 VPWR.n2 VPWR.t27 381.443
R90 VPWR.n324 VPWR.t28 381.443
R91 VPWR.n0 VPWR.t72 381.443
R92 VPWR.n726 VPWR.t73 381.443
R93 VPWR.n421 VPWR.t140 381.443
R94 VPWR.n18 VPWR.t83 380.193
R95 VPWR.n21 VPWR.t90 380.193
R96 VPWR.n499 VPWR.t44 380.193
R97 VPWR.n502 VPWR.t52 380.193
R98 VPWR.n78 VPWR.t55 380.193
R99 VPWR.n81 VPWR.t97 380.193
R100 VPWR.n573 VPWR.t29 380.193
R101 VPWR.n576 VPWR.t7 380.193
R102 VPWR.n183 VPWR.t158 380.193
R103 VPWR.n186 VPWR.t142 380.193
R104 VPWR.n606 VPWR.t202 380.193
R105 VPWR.n609 VPWR.t21 380.193
R106 VPWR.t133 VPWR 369.938
R107 VPWR VPWR.t153 366.978
R108 VPWR VPWR.t57 357.51
R109 VPWR.n77 VPWR.t188 344.06
R110 VPWR.n192 VPWR.t209 344.06
R111 VPWR.n261 VPWR.t42 344.06
R112 VPWR.n192 VPWR.t61 344.06
R113 VPWR.n230 VPWR.t77 344.06
R114 VPWR.n28 VPWR.t13 340.243
R115 VPWR.n29 VPWR.t120 338.488
R116 VPWR VPWR.t54 334.012
R117 VPWR VPWR.t26 322.587
R118 VPWR.n316 VPWR 322.587
R119 VPWR.t138 VPWR 322.587
R120 VPWR.n113 VPWR.n66 322.329
R121 VPWR.n36 VPWR.n35 320.976
R122 VPWR.n38 VPWR.n37 320.976
R123 VPWR.n33 VPWR.n16 320.976
R124 VPWR.n338 VPWR.n321 315.406
R125 VPWR.n417 VPWR.n286 312.053
R126 VPWR.n308 VPWR.n307 312.053
R127 VPWR.n169 VPWR.n168 312.005
R128 VPWR.n270 VPWR.n269 311.892
R129 VPWR.n173 VPWR.n172 311.659
R130 VPWR.n173 VPWR.n171 311.659
R131 VPWR.n215 VPWR.n214 311.519
R132 VPWR.n636 VPWR.n266 310.5
R133 VPWR.n705 VPWR.n34 308.151
R134 VPWR.n105 VPWR.n69 308.151
R135 VPWR.n273 VPWR.n272 308.151
R136 VPWR.n244 VPWR.n158 308.149
R137 VPWR.n451 VPWR.t222 306.735
R138 VPWR.n451 VPWR.t236 306.735
R139 VPWR.n489 VPWR.t224 306.735
R140 VPWR.n489 VPWR.t241 306.735
R141 VPWR.n667 VPWR.t229 306.735
R142 VPWR.n107 VPWR.t218 306.735
R143 VPWR.n142 VPWR.t237 306.735
R144 VPWR.n556 VPWR.t231 306.735
R145 VPWR.n156 VPWR.t235 306.735
R146 VPWR.n380 VPWR.t245 306.735
R147 VPWR.t199 VPWR.t115 298.764
R148 VPWR.t31 VPWR.t179 298.764
R149 VPWR.t111 VPWR.t133 290.031
R150 VPWR.t211 VPWR.t160 281.154
R151 VPWR.t151 VPWR.t99 281.154
R152 VPWR VPWR.t43 280.3
R153 VPWR VPWR.t6 280.3
R154 VPWR VPWR.t20 278.623
R155 VPWR VPWR.t204 260.159
R156 VPWR.n287 VPWR.t154 249.363
R157 VPWR.n364 VPWR.t163 249.363
R158 VPWR.t160 VPWR.t162 248.599
R159 VPWR.t153 VPWR.t151 248.599
R160 VPWR.n697 VPWR.t175 246.817
R161 VPWR.n19 VPWR.t240 245.667
R162 VPWR.n22 VPWR.t223 245.667
R163 VPWR.n500 VPWR.t244 245.667
R164 VPWR.n503 VPWR.t227 245.667
R165 VPWR.n79 VPWR.t230 245.667
R166 VPWR.n82 VPWR.t247 245.667
R167 VPWR.n574 VPWR.t233 245.667
R168 VPWR.n577 VPWR.t220 245.667
R169 VPWR.n184 VPWR.t246 245.667
R170 VPWR.n187 VPWR.t238 245.667
R171 VPWR.n607 VPWR.t219 245.667
R172 VPWR.n610 VPWR.t242 245.667
R173 VPWR.n420 VPWR.t234 242.282
R174 VPWR.n322 VPWR.t228 242.282
R175 VPWR.n727 VPWR.t232 242.282
R176 VPWR.t71 VPWR 221.964
R177 VPWR.n316 VPWR 219.004
R178 VPWR.n41 VPWR.t226 215.827
R179 VPWR.n695 VPWR.t221 214.929
R180 VPWR.n166 VPWR.n165 213.119
R181 VPWR.n349 VPWR.n316 213.119
R182 VPWR.t135 VPWR.t111 213.084
R183 VPWR.n370 VPWR.t243 210.964
R184 VPWR.n689 VPWR.n45 210.55
R185 VPWR.t88 VPWR 209.806
R186 VPWR.n121 VPWR.n63 209.368
R187 VPWR.t23 VPWR 203.093
R188 VPWR VPWR.t215 203.093
R189 VPWR VPWR.t49 203.093
R190 VPWR VPWR.t144 203.093
R191 VPWR.t99 VPWR 192.369
R192 VPWR VPWR.t166 189.409
R193 VPWR.t43 VPWR 182.952
R194 VPWR.n63 VPWR 182.952
R195 VPWR.t6 VPWR 182.952
R196 VPWR.t20 VPWR 182.952
R197 VPWR.t172 VPWR.t129 181.273
R198 VPWR.n45 VPWR 179.595
R199 VPWR VPWR.t178 177.916
R200 VPWR VPWR.t109 169.524
R201 VPWR.t0 VPWR.t168 164.488
R202 VPWR.t2 VPWR.t113 164.488
R203 VPWR.t33 VPWR.t193 161.131
R204 VPWR.t4 VPWR.t66 161.131
R205 VPWR.t74 VPWR.t197 161.131
R206 VPWR.n563 VPWR.n562 159.476
R207 VPWR.n252 VPWR.n251 159.476
R208 VPWR.t115 VPWR.t0 147.703
R209 VPWR.t179 VPWR.t2 147.703
R210 VPWR.t189 VPWR.t187 144.346
R211 VPWR.t191 VPWR.t189 144.346
R212 VPWR.t193 VPWR.t191 144.346
R213 VPWR.t62 VPWR.t60 144.346
R214 VPWR.t64 VPWR.t62 144.346
R215 VPWR.t66 VPWR.t64 144.346
R216 VPWR.t76 VPWR.t78 144.346
R217 VPWR.t78 VPWR.t80 144.346
R218 VPWR.t80 VPWR.t74 144.346
R219 VPWR.t174 VPWR.t181 140.989
R220 VPWR.t109 VPWR.t172 140.989
R221 VPWR.t107 VPWR.t121 140.989
R222 VPWR.t171 VPWR.t186 140.989
R223 VPWR.t186 VPWR.t170 140.989
R224 VPWR.t170 VPWR.t185 140.989
R225 VPWR.t37 VPWR.t127 139.311
R226 VPWR.t39 VPWR.t125 135.954
R227 VPWR.n627 VPWR.t239 129.344
R228 VPWR.t82 VPWR 125.883
R229 VPWR.t54 VPWR 125.883
R230 VPWR.n63 VPWR 125.883
R231 VPWR.t141 VPWR 125.883
R232 VPWR.n60 VPWR.t225 124.891
R233 VPWR.n66 VPWR.t173 116.341
R234 VPWR VPWR.t33 110.778
R235 VPWR VPWR.t4 110.778
R236 VPWR.t197 VPWR 110.778
R237 VPWR.t136 VPWR 110.778
R238 VPWR.t168 VPWR 109.1
R239 VPWR.t113 VPWR 109.1
R240 VPWR VPWR.t174 107.421
R241 VPWR.t147 VPWR 105.743
R242 VPWR.t131 VPWR.t88 100.707
R243 VPWR.t195 VPWR.t123 99.0288
R244 VPWR.t101 VPWR.t176 99.0288
R245 VPWR.t178 VPWR.t201 99.0288
R246 VPWR.n570 VPWR.t1 96.1553
R247 VPWR.n214 VPWR.t177 96.1553
R248 VPWR.n168 VPWR.t102 96.1553
R249 VPWR.n153 VPWR.t3 96.1553
R250 VPWR.n321 VPWR.t112 96.1553
R251 VPWR VPWR.t211 91.745
R252 VPWR.t41 VPWR 88.9581
R253 VPWR.n562 VPWR.t116 86.7743
R254 VPWR.n251 VPWR.t180 86.7743
R255 VPWR.t185 VPWR.t46 83.9228
R256 VPWR.n165 VPWR.t105 80.5659
R257 VPWR.t18 VPWR.t117 78.8874
R258 VPWR VPWR.t164 78.8874
R259 VPWR.n45 VPWR.t9 77.209
R260 VPWR.t129 VPWR.t23 77.209
R261 VPWR.t16 VPWR.t103 75.5305
R262 VPWR.t119 VPWR.t12 72.1736
R263 VPWR.t14 VPWR.t119 72.1736
R264 VPWR.t164 VPWR 72.1736
R265 VPWR.t187 VPWR 70.4952
R266 VPWR VPWR.t76 70.4952
R267 VPWR.t103 VPWR.t14 68.8168
R268 VPWR VPWR.t183 68.8168
R269 VPWR.n563 VPWR.t200 66.8398
R270 VPWR.n252 VPWR.t32 66.8398
R271 VPWR.t117 VPWR.t16 65.4599
R272 VPWR VPWR.t41 65.4599
R273 VPWR.t176 VPWR.t131 63.7814
R274 VPWR.n570 VPWR.t169 63.3219
R275 VPWR.n153 VPWR.t114 63.3219
R276 VPWR.t123 VPWR.t18 62.103
R277 VPWR.t181 VPWR 62.103
R278 VPWR.n286 VPWR.t100 55.4067
R279 VPWR.n307 VPWR.t212 55.4067
R280 VPWR VPWR.t35 55.3892
R281 VPWR.n61 VPWR.n60 50.7764
R282 VPWR.t204 VPWR 50.3539
R283 VPWR.t9 VPWR 48.6754
R284 VPWR.t105 VPWR 45.3185
R285 VPWR.t183 VPWR.t195 41.9616
R286 VPWR.n34 VPWR.t19 37.4305
R287 VPWR.n69 VPWR.t194 37.4305
R288 VPWR.n171 VPWR.t67 37.4305
R289 VPWR.n172 VPWR.t208 37.4305
R290 VPWR.n158 VPWR.t75 37.4305
R291 VPWR.n272 VPWR.t40 37.4305
R292 VPWR.n701 VPWR.n700 34.6358
R293 VPWR.n31 VPWR.n30 34.6358
R294 VPWR.n213 VPWR.n212 34.6358
R295 VPWR.n216 VPWR.n213 34.6358
R296 VPWR.n220 VPWR.n219 34.6358
R297 VPWR.n221 VPWR.n220 34.6358
R298 VPWR.n632 VPWR.n631 34.6358
R299 VPWR.n348 VPWR.n317 34.6358
R300 VPWR.n342 VPWR.n319 34.6358
R301 VPWR.n343 VPWR.n342 34.6358
R302 VPWR.n286 VPWR.t152 34.0906
R303 VPWR.n307 VPWR.t161 34.0906
R304 VPWR.n706 VPWR.n705 32.377
R305 VPWR.n66 VPWR.t130 28.4453
R306 VPWR.n34 VPWR.t196 27.5805
R307 VPWR.n17 VPWR.t15 27.5805
R308 VPWR.n17 VPWR.t17 27.5805
R309 VPWR.n69 VPWR.t34 27.5805
R310 VPWR.n70 VPWR.t190 27.5805
R311 VPWR.n70 VPWR.t192 27.5805
R312 VPWR.n194 VPWR.t63 27.5805
R313 VPWR.n194 VPWR.t65 27.5805
R314 VPWR.n195 VPWR.t210 27.5805
R315 VPWR.n195 VPWR.t207 27.5805
R316 VPWR.n171 VPWR.t5 27.5805
R317 VPWR.n172 VPWR.t150 27.5805
R318 VPWR.n159 VPWR.t79 27.5805
R319 VPWR.n159 VPWR.t81 27.5805
R320 VPWR.n158 VPWR.t198 27.5805
R321 VPWR.n268 VPWR.t36 27.5805
R322 VPWR.n268 VPWR.t38 27.5805
R323 VPWR.n272 VPWR.t137 27.5805
R324 VPWR.n165 VPWR 26.8556
R325 VPWR.n214 VPWR.t89 26.5955
R326 VPWR.n321 VPWR.t134 26.5955
R327 VPWR.n35 VPWR.t124 26.5955
R328 VPWR.n35 VPWR.t184 26.5955
R329 VPWR.n37 VPWR.t165 26.5955
R330 VPWR.n37 VPWR.t182 26.5955
R331 VPWR.n16 VPWR.t104 26.5955
R332 VPWR.n16 VPWR.t118 26.5955
R333 VPWR.n266 VPWR.t108 26.5955
R334 VPWR.n266 VPWR.t122 26.5955
R335 VPWR.n269 VPWR.t128 26.5955
R336 VPWR.n269 VPWR.t126 26.5955
R337 VPWR.n635 VPWR.n270 26.3534
R338 VPWR.n124 VPWR.n123 26.3341
R339 VPWR.n344 VPWR.n343 25.977
R340 VPWR.n168 VPWR.t132 25.6105
R341 VPWR.n197 VPWR.n193 25.6005
R342 VPWR.n416 VPWR.n287 25.6005
R343 VPWR.n364 VPWR.n363 25.6005
R344 VPWR.n212 VPWR.n173 25.224
R345 VPWR.n338 VPWR.n337 25.224
R346 VPWR.n631 VPWR.n630 25.1912
R347 VPWR.n426 VPWR.n425 25.1912
R348 VPWR.n368 VPWR.n305 25.1912
R349 VPWR.n337 VPWR.n325 25.1912
R350 VPWR.t125 VPWR.t136 25.1772
R351 VPWR.n701 VPWR.n36 24.8476
R352 VPWR.n426 VPWR.n417 24.8476
R353 VPWR.n350 VPWR.n308 24.8476
R354 VPWR.n197 VPWR.n196 24.4711
R355 VPWR.n364 VPWR.n305 24.0946
R356 VPWR.n344 VPWR.n317 24.0946
R357 VPWR.n27 VPWR.n24 23.7181
R358 VPWR.n221 VPWR.n166 23.7181
R359 VPWR.n350 VPWR.n349 23.7181
R360 VPWR.n349 VPWR.n348 23.7181
R361 VPWR.n637 VPWR.n636 22.9652
R362 VPWR.n338 VPWR.n319 22.9652
R363 VPWR.t201 VPWR.t101 21.8203
R364 VPWR.n215 VPWR.n169 21.4593
R365 VPWR.n636 VPWR.n635 21.4593
R366 VPWR.n196 VPWR.n173 20.7064
R367 VPWR.n135 VPWR.n61 20.0749
R368 VPWR.n645 VPWR.n261 20.0094
R369 VPWR.n697 VPWR.n38 19.9534
R370 VPWR.n193 VPWR.n192 19.9534
R371 VPWR.n637 VPWR.n261 19.9534
R372 VPWR.n417 VPWR.n416 19.577
R373 VPWR.n363 VPWR.n308 19.577
R374 VPWR.n706 VPWR.n33 18.824
R375 VPWR.n377 VPWR.n304 17.612
R376 VPWR.n84 VPWR.n77 16.9417
R377 VPWR.n192 VPWR.n189 16.9417
R378 VPWR.n230 VPWR.n166 16.9417
R379 VPWR.n482 VPWR.n481 16.6847
R380 VPWR.n404 VPWR.n287 16.2447
R381 VPWR.n581 VPWR.n580 15.8683
R382 VPWR.n30 VPWR.n29 15.8123
R383 VPWR.n725 VPWR.n724 15.7465
R384 VPWR.n33 VPWR.n32 15.0593
R385 VPWR.n689 VPWR.n688 14.9
R386 VPWR.n29 VPWR.n28 14.6829
R387 VPWR.n507 VPWR.n506 14.5851
R388 VPWR.n614 VPWR.n613 14.2735
R389 VPWR.n92 VPWR.n77 12.3742
R390 VPWR.n231 VPWR.n230 12.3742
R391 VPWR.n219 VPWR.n169 12.0476
R392 VPWR.n704 VPWR.n36 9.78874
R393 VPWR.n108 VPWR.n67 9.73273
R394 VPWR.n112 VPWR.n67 9.73273
R395 VPWR.n116 VPWR.n114 9.73273
R396 VPWR.n121 VPWR.n64 9.73273
R397 VPWR.n592 VPWR.n569 9.73273
R398 VPWR.n249 VPWR.n248 9.73273
R399 VPWR.n259 VPWR.n258 9.73273
R400 VPWR.n383 VPWR.n379 9.73273
R401 VPWR.n383 VPWR.n382 9.73273
R402 VPWR.n395 VPWR.n293 9.73273
R403 VPWR.n396 VPWR.n395 9.73273
R404 VPWR.n397 VPWR.n396 9.73273
R405 VPWR.n397 VPWR.n291 9.73273
R406 VPWR.n401 VPWR.n291 9.73273
R407 VPWR.n402 VPWR.n401 9.73273
R408 VPWR VPWR.n0 9.6274
R409 VPWR.n421 VPWR.n419 9.60526
R410 VPWR.n104 VPWR.n71 9.52116
R411 VPWR.n591 VPWR.n590 9.52116
R412 VPWR.n243 VPWR.n242 9.52116
R413 VPWR.n647 VPWR.n260 9.52116
R414 VPWR.n124 VPWR.n122 9.49016
R415 VPWR.n27 VPWR.n26 9.3005
R416 VPWR.n30 VPWR.n12 9.3005
R417 VPWR.n31 VPWR.n13 9.3005
R418 VPWR.n707 VPWR.n706 9.3005
R419 VPWR.n704 VPWR.n703 9.3005
R420 VPWR.n702 VPWR.n701 9.3005
R421 VPWR.n700 VPWR.n699 9.3005
R422 VPWR.n690 VPWR.n689 9.3005
R423 VPWR.n689 VPWR.n44 9.3005
R424 VPWR.n688 VPWR.n687 9.3005
R425 VPWR.n453 VPWR.n48 9.3005
R426 VPWR.n454 VPWR.n452 9.3005
R427 VPWR.n456 VPWR.n455 9.3005
R428 VPWR.n458 VPWR.n457 9.3005
R429 VPWR.n459 VPWR.n450 9.3005
R430 VPWR.n461 VPWR.n460 9.3005
R431 VPWR.n462 VPWR.n449 9.3005
R432 VPWR.n465 VPWR.n464 9.3005
R433 VPWR.n466 VPWR.n448 9.3005
R434 VPWR.n468 VPWR.n467 9.3005
R435 VPWR.n481 VPWR.n480 9.3005
R436 VPWR.n482 VPWR.n441 9.3005
R437 VPWR.n485 VPWR.n484 9.3005
R438 VPWR.n486 VPWR.n440 9.3005
R439 VPWR.n488 VPWR.n487 9.3005
R440 VPWR.n490 VPWR.n439 9.3005
R441 VPWR.n492 VPWR.n491 9.3005
R442 VPWR.n493 VPWR.n438 9.3005
R443 VPWR.n495 VPWR.n494 9.3005
R444 VPWR.n496 VPWR.n436 9.3005
R445 VPWR.n518 VPWR.n517 9.3005
R446 VPWR.n516 VPWR.n515 9.3005
R447 VPWR.n508 VPWR.n507 9.3005
R448 VPWR.n86 VPWR.n77 9.3005
R449 VPWR.n92 VPWR.n91 9.3005
R450 VPWR.n95 VPWR.n94 9.3005
R451 VPWR.n104 VPWR.n103 9.3005
R452 VPWR.n106 VPWR.n68 9.3005
R453 VPWR.n109 VPWR.n108 9.3005
R454 VPWR.n110 VPWR.n67 9.3005
R455 VPWR.n112 VPWR.n111 9.3005
R456 VPWR.n114 VPWR.n65 9.3005
R457 VPWR.n117 VPWR.n116 9.3005
R458 VPWR.n118 VPWR.n64 9.3005
R459 VPWR.n121 VPWR.n120 9.3005
R460 VPWR.n125 VPWR.n124 9.3005
R461 VPWR.n135 VPWR.n134 9.3005
R462 VPWR.n138 VPWR.n58 9.3005
R463 VPWR.n670 VPWR.n669 9.3005
R464 VPWR.n668 VPWR.n59 9.3005
R465 VPWR.n665 VPWR.n664 9.3005
R466 VPWR.n663 VPWR.n139 9.3005
R467 VPWR.n662 VPWR.n661 9.3005
R468 VPWR.n660 VPWR.n140 9.3005
R469 VPWR.n659 VPWR.n658 9.3005
R470 VPWR.n538 VPWR.n143 9.3005
R471 VPWR.n540 VPWR.n539 9.3005
R472 VPWR.n550 VPWR.n549 9.3005
R473 VPWR.n552 VPWR.n551 9.3005
R474 VPWR.n554 VPWR.n553 9.3005
R475 VPWR.n555 VPWR.n533 9.3005
R476 VPWR.n558 VPWR.n557 9.3005
R477 VPWR.n560 VPWR.n559 9.3005
R478 VPWR.n561 VPWR.n531 9.3005
R479 VPWR.n566 VPWR.n565 9.3005
R480 VPWR.n568 VPWR.n567 9.3005
R481 VPWR.n569 VPWR.n528 9.3005
R482 VPWR.n593 VPWR.n592 9.3005
R483 VPWR.n590 VPWR.n589 9.3005
R484 VPWR.n582 VPWR.n581 9.3005
R485 VPWR.n192 VPWR.n191 9.3005
R486 VPWR.n193 VPWR.n181 9.3005
R487 VPWR.n198 VPWR.n197 9.3005
R488 VPWR.n196 VPWR.n174 9.3005
R489 VPWR.n210 VPWR.n173 9.3005
R490 VPWR.n212 VPWR.n211 9.3005
R491 VPWR.n213 VPWR.n170 9.3005
R492 VPWR.n217 VPWR.n216 9.3005
R493 VPWR.n219 VPWR.n218 9.3005
R494 VPWR.n220 VPWR.n167 9.3005
R495 VPWR.n222 VPWR.n221 9.3005
R496 VPWR.n223 VPWR.n166 9.3005
R497 VPWR.n230 VPWR.n229 9.3005
R498 VPWR.n232 VPWR.n231 9.3005
R499 VPWR.n241 VPWR.n240 9.3005
R500 VPWR.n243 VPWR.n157 9.3005
R501 VPWR.n246 VPWR.n245 9.3005
R502 VPWR.n248 VPWR.n247 9.3005
R503 VPWR.n249 VPWR.n155 9.3005
R504 VPWR.n255 VPWR.n254 9.3005
R505 VPWR.n256 VPWR.n154 9.3005
R506 VPWR.n258 VPWR.n257 9.3005
R507 VPWR.n259 VPWR.n152 9.3005
R508 VPWR.n648 VPWR.n647 9.3005
R509 VPWR.n645 VPWR.n644 9.3005
R510 VPWR.n639 VPWR.n261 9.3005
R511 VPWR.n638 VPWR.n637 9.3005
R512 VPWR.n636 VPWR.n267 9.3005
R513 VPWR.n635 VPWR.n634 9.3005
R514 VPWR.n633 VPWR.n632 9.3005
R515 VPWR.n631 VPWR.n271 9.3005
R516 VPWR.n630 VPWR.n629 9.3005
R517 VPWR.n628 VPWR.n627 9.3005
R518 VPWR.n626 VPWR.n625 9.3005
R519 VPWR.n277 VPWR.n276 9.3005
R520 VPWR.n604 VPWR.n603 9.3005
R521 VPWR.n615 VPWR.n614 9.3005
R522 VPWR.n729 VPWR.n728 9.3005
R523 VPWR.n725 VPWR.n1 9.3005
R524 VPWR.n724 VPWR.n723 9.3005
R525 VPWR.n323 VPWR.n3 9.3005
R526 VPWR.n328 VPWR.n325 9.3005
R527 VPWR.n337 VPWR.n336 9.3005
R528 VPWR.n339 VPWR.n338 9.3005
R529 VPWR.n340 VPWR.n319 9.3005
R530 VPWR.n342 VPWR.n341 9.3005
R531 VPWR.n343 VPWR.n318 9.3005
R532 VPWR.n345 VPWR.n344 9.3005
R533 VPWR.n346 VPWR.n317 9.3005
R534 VPWR.n348 VPWR.n347 9.3005
R535 VPWR.n349 VPWR.n315 9.3005
R536 VPWR.n351 VPWR.n350 9.3005
R537 VPWR.n309 VPWR.n308 9.3005
R538 VPWR.n363 VPWR.n362 9.3005
R539 VPWR.n365 VPWR.n364 9.3005
R540 VPWR.n366 VPWR.n305 9.3005
R541 VPWR.n368 VPWR.n367 9.3005
R542 VPWR.n371 VPWR 9.3005
R543 VPWR.n374 VPWR.n373 9.3005
R544 VPWR.n375 VPWR.n304 9.3005
R545 VPWR.n377 VPWR.n376 9.3005
R546 VPWR.n379 VPWR.n300 9.3005
R547 VPWR.n384 VPWR.n383 9.3005
R548 VPWR.n382 VPWR.n381 9.3005
R549 VPWR.n393 VPWR.n293 9.3005
R550 VPWR.n395 VPWR.n394 9.3005
R551 VPWR.n396 VPWR.n292 9.3005
R552 VPWR.n398 VPWR.n397 9.3005
R553 VPWR.n399 VPWR.n291 9.3005
R554 VPWR.n401 VPWR.n400 9.3005
R555 VPWR.n402 VPWR.n290 9.3005
R556 VPWR.n405 VPWR.n404 9.3005
R557 VPWR.n406 VPWR.n287 9.3005
R558 VPWR.n416 VPWR.n415 9.3005
R559 VPWR.n417 VPWR.n285 9.3005
R560 VPWR.n427 VPWR.n426 9.3005
R561 VPWR.n425 VPWR.n424 9.3005
R562 VPWR.n423 VPWR.n422 9.3005
R563 VPWR.n94 VPWR.n93 9.09802
R564 VPWR.n105 VPWR.n104 9.09802
R565 VPWR.n590 VPWR.n571 9.09802
R566 VPWR.n241 VPWR.n160 9.09802
R567 VPWR.n244 VPWR.n243 9.09802
R568 VPWR.n647 VPWR.n646 9.09802
R569 VPWR.n379 VPWR.n378 9.09802
R570 VPWR.n403 VPWR.n402 9.09802
R571 VPWR.n123 VPWR.n61 8.9761
R572 VPWR.n565 VPWR.n561 8.80773
R573 VPWR.n254 VPWR.n249 8.80773
R574 VPWR.n569 VPWR.n568 8.57648
R575 VPWR.n258 VPWR.n154 8.57648
R576 VPWR.n561 VPWR.n560 8.44958
R577 VPWR.n693 VPWR.n692 7.93422
R578 VPWR.n551 VPWR.n550 7.21067
R579 VPWR.n122 VPWR.n121 6.66496
R580 VPWR.n665 VPWR.n139 6.52104
R581 VPWR.n692 VPWR.n39 6.48583
R582 VPWR.n689 VPWR.n43 6.46951
R583 VPWR.n273 VPWR.n270 6.02403
R584 VPWR.n42 VPWR.n41 5.8885
R585 VPWR.n454 VPWR.n453 5.66204
R586 VPWR.n455 VPWR.n454 5.66204
R587 VPWR.n459 VPWR.n458 5.66204
R588 VPWR.n460 VPWR.n459 5.66204
R589 VPWR.n460 VPWR.n449 5.66204
R590 VPWR.n465 VPWR.n449 5.66204
R591 VPWR.n466 VPWR.n465 5.66204
R592 VPWR.n467 VPWR.n466 5.66204
R593 VPWR.n484 VPWR.n440 5.66204
R594 VPWR.n488 VPWR.n440 5.66204
R595 VPWR.n491 VPWR.n490 5.66204
R596 VPWR.n491 VPWR.n438 5.66204
R597 VPWR.n495 VPWR.n438 5.66204
R598 VPWR.n496 VPWR.n495 5.66204
R599 VPWR.n517 VPWR.n496 5.66204
R600 VPWR.n517 VPWR.n516 5.66204
R601 VPWR.n661 VPWR.n660 5.66204
R602 VPWR.n660 VPWR.n659 5.66204
R603 VPWR.n539 VPWR.n538 5.66204
R604 VPWR.n555 VPWR.n554 5.66204
R605 VPWR.n557 VPWR.n555 5.66204
R606 VPWR.n116 VPWR.n115 5.60711
R607 VPWR.n453 VPWR.n46 5.29281
R608 VPWR.n467 VPWR.n442 5.29281
R609 VPWR.n484 VPWR.n483 5.29281
R610 VPWR.n516 VPWR.n497 5.29281
R611 VPWR.n661 VPWR.n141 5.29281
R612 VPWR.n539 VPWR.n536 5.29281
R613 VPWR.n554 VPWR.n534 5.29281
R614 VPWR.n114 VPWR.n113 5.28976
R615 VPWR.n697 VPWR.n696 5.28746
R616 VPWR.n107 VPWR.n106 5.18397
R617 VPWR.n245 VPWR.n156 5.18397
R618 VPWR.n382 VPWR.n380 5.18397
R619 VPWR.t127 VPWR.t39 5.03584
R620 VPWR VPWR.t171 5.03584
R621 VPWR.n695 VPWR.n694 4.8005
R622 VPWR.n627 VPWR.n626 4.67352
R623 VPWR.n626 VPWR.n276 4.67352
R624 VPWR.n604 VPWR.n276 4.67352
R625 VPWR.n373 VPWR.n371 4.67352
R626 VPWR.n698 VPWR.n697 4.62124
R627 VPWR.n692 VPWR.n691 4.62124
R628 VPWR.n108 VPWR.n107 4.54926
R629 VPWR.n248 VPWR.n156 4.54926
R630 VPWR.n380 VPWR.n293 4.54926
R631 VPWR.n722 VPWR.n721 4.51401
R632 VPWR.n333 VPWR.n320 4.51401
R633 VPWR.n354 VPWR.n312 4.51401
R634 VPWR.n359 VPWR.n306 4.51401
R635 VPWR.n387 VPWR.n298 4.51401
R636 VPWR.n392 VPWR.n391 4.51401
R637 VPWR.n657 VPWR.n656 4.51401
R638 VPWR.n546 VPWR.n535 4.51401
R639 VPWR.n651 VPWR.n150 4.51401
R640 VPWR.n641 VPWR.n640 4.51401
R641 VPWR.n463 VPWR.n447 4.51401
R642 VPWR.n477 VPWR.n445 4.51401
R643 VPWR.n716 VPWR.n10 4.51401
R644 VPWR.n15 VPWR.n14 4.51401
R645 VPWR.n521 VPWR.n434 4.51401
R646 VPWR.n514 VPWR.n513 4.51401
R647 VPWR.n680 VPWR.n40 4.51401
R648 VPWR.n684 VPWR.n50 4.51401
R649 VPWR.n226 VPWR.n224 4.51401
R650 VPWR.n239 VPWR.n238 4.51401
R651 VPWR.n119 VPWR.n62 4.51401
R652 VPWR.n672 VPWR.n671 4.51401
R653 VPWR.n596 VPWR.n526 4.51401
R654 VPWR.n588 VPWR.n587 4.51401
R655 VPWR.n90 VPWR.n89 4.51401
R656 VPWR.n102 VPWR.n101 4.51401
R657 VPWR.n204 VPWR.n179 4.51401
R658 VPWR.n209 VPWR.n208 4.51401
R659 VPWR.n278 VPWR.n275 4.51401
R660 VPWR.n617 VPWR.n616 4.51401
R661 VPWR.n408 VPWR.n407 4.51401
R662 VPWR.n429 VPWR.n428 4.51401
R663 VPWR.n512 VPWR.n498 4.5005
R664 VPWR.n715 VPWR.n714 4.5005
R665 VPWR.n713 VPWR.n712 4.5005
R666 VPWR.n709 VPWR.n708 4.5005
R667 VPWR.n470 VPWR.n469 4.5005
R668 VPWR.n471 VPWR.n443 4.5005
R669 VPWR.n479 VPWR.n478 4.5005
R670 VPWR.n520 VPWR.n519 4.5005
R671 VPWR.n509 VPWR.n437 4.5005
R672 VPWR.n679 VPWR.n678 4.5005
R673 VPWR.n676 VPWR.n47 4.5005
R674 VPWR.n686 VPWR.n685 4.5005
R675 VPWR.n586 VPWR.n572 4.5005
R676 VPWR.n127 VPWR.n126 4.5005
R677 VPWR.n132 VPWR.n131 4.5005
R678 VPWR.n133 VPWR.n57 4.5005
R679 VPWR.n537 VPWR.n144 4.5005
R680 VPWR.n543 VPWR.n541 4.5005
R681 VPWR.n548 VPWR.n547 4.5005
R682 VPWR.n595 VPWR.n594 4.5005
R683 VPWR.n583 VPWR.n529 4.5005
R684 VPWR.n87 VPWR.n76 4.5005
R685 VPWR.n97 VPWR.n96 4.5005
R686 VPWR.n73 VPWR.n72 4.5005
R687 VPWR.n203 VPWR.n202 4.5005
R688 VPWR.n201 VPWR.n200 4.5005
R689 VPWR.n182 VPWR.n175 4.5005
R690 VPWR.n228 VPWR.n227 4.5005
R691 VPWR.n234 VPWR.n233 4.5005
R692 VPWR.n162 VPWR.n161 4.5005
R693 VPWR.n650 VPWR.n649 4.5005
R694 VPWR.n263 VPWR.n262 4.5005
R695 VPWR.n643 VPWR.n642 4.5005
R696 VPWR.n602 VPWR.n600 4.5005
R697 VPWR.n624 VPWR.n623 4.5005
R698 VPWR.n601 VPWR.n279 4.5005
R699 VPWR.n289 VPWR.n284 4.5005
R700 VPWR.n327 VPWR.n4 4.5005
R701 VPWR.n330 VPWR.n329 4.5005
R702 VPWR.n335 VPWR.n334 4.5005
R703 VPWR.n353 VPWR.n352 4.5005
R704 VPWR.n314 VPWR.n313 4.5005
R705 VPWR.n361 VPWR.n360 4.5005
R706 VPWR.n386 VPWR.n385 4.5005
R707 VPWR.n303 VPWR.n302 4.5005
R708 VPWR.n295 VPWR.n294 4.5005
R709 VPWR.n409 VPWR.n288 4.5005
R710 VPWR.n414 VPWR.n413 4.5005
R711 VPWR.n113 VPWR.n112 4.44348
R712 VPWR.n627 VPWR.n274 4.36875
R713 VPWR.n605 VPWR.n604 4.36875
R714 VPWR.n422 VPWR.n421 4.36875
R715 VPWR.n373 VPWR.n372 4.36875
R716 VPWR.n324 VPWR.n323 4.36875
R717 VPWR.n728 VPWR.n0 4.36875
R718 VPWR.n137 VPWR.n60 4.31787
R719 VPWR.n28 VPWR.n27 4.14168
R720 VPWR.n115 VPWR.n64 4.12612
R721 VPWR.n564 VPWR.n530 4.04887
R722 VPWR.n253 VPWR.n250 4.04887
R723 VPWR.n24 VPWR.n20 4.02033
R724 VPWR.n24 VPWR.n23 4.02033
R725 VPWR.n506 VPWR.n501 4.02033
R726 VPWR.n506 VPWR.n504 4.02033
R727 VPWR.n84 VPWR.n80 4.02033
R728 VPWR.n84 VPWR.n83 4.02033
R729 VPWR.n580 VPWR.n575 4.02033
R730 VPWR.n580 VPWR.n578 4.02033
R731 VPWR.n189 VPWR.n185 4.02033
R732 VPWR.n189 VPWR.n188 4.02033
R733 VPWR.n613 VPWR.n608 4.02033
R734 VPWR.n613 VPWR.n611 4.02033
R735 VPWR.n700 VPWR.n38 3.76521
R736 VPWR.n422 VPWR.n420 3.50526
R737 VPWR.n323 VPWR.n322 3.50526
R738 VPWR.n728 VPWR.n727 3.50526
R739 VPWR.n669 VPWR.n138 3.47425
R740 VPWR.n669 VPWR.n668 3.47425
R741 VPWR.n333 VPWR.n6 3.43925
R742 VPWR.n721 VPWR.n720 3.43925
R743 VPWR.n359 VPWR.n358 3.43925
R744 VPWR.n355 VPWR.n354 3.43925
R745 VPWR.n391 VPWR.n390 3.43925
R746 VPWR.n388 VPWR.n387 3.43925
R747 VPWR.n546 VPWR.n147 3.43925
R748 VPWR.n656 VPWR.n655 3.43925
R749 VPWR.n641 VPWR.n148 3.43925
R750 VPWR.n652 VPWR.n651 3.43925
R751 VPWR.n14 VPWR.n7 3.43925
R752 VPWR.n717 VPWR.n716 3.43925
R753 VPWR.n513 VPWR.n432 3.43925
R754 VPWR.n522 VPWR.n521 3.43925
R755 VPWR.n684 VPWR.n683 3.43925
R756 VPWR.n681 VPWR.n680 3.43925
R757 VPWR.n238 VPWR.n237 3.43925
R758 VPWR.n226 VPWR.n225 3.43925
R759 VPWR.n587 VPWR.n524 3.43925
R760 VPWR.n597 VPWR.n596 3.43925
R761 VPWR.n101 VPWR.n100 3.43925
R762 VPWR.n89 VPWR.n88 3.43925
R763 VPWR.n618 VPWR.n617 3.43925
R764 VPWR.n620 VPWR.n278 3.43925
R765 VPWR.n326 VPWR.n5 3.4105
R766 VPWR.n332 VPWR.n331 3.4105
R767 VPWR.n356 VPWR.n311 3.4105
R768 VPWR.n357 VPWR.n310 3.4105
R769 VPWR.n299 VPWR.n297 3.4105
R770 VPWR.n301 VPWR.n296 3.4105
R771 VPWR.n542 VPWR.n145 3.4105
R772 VPWR.n545 VPWR.n544 3.4105
R773 VPWR.n151 VPWR.n149 3.4105
R774 VPWR.n265 VPWR.n264 3.4105
R775 VPWR.n476 VPWR.n146 3.4105
R776 VPWR.n446 VPWR.n146 3.4105
R777 VPWR.n477 VPWR.n476 3.4105
R778 VPWR.n447 VPWR.n446 3.4105
R779 VPWR.n473 VPWR.n472 3.4105
R780 VPWR.n475 VPWR.n444 3.4105
R781 VPWR.n11 VPWR.n9 3.4105
R782 VPWR.n711 VPWR.n710 3.4105
R783 VPWR.n435 VPWR.n433 3.4105
R784 VPWR.n511 VPWR.n510 3.4105
R785 VPWR.n677 VPWR.n675 3.4105
R786 VPWR.n51 VPWR.n49 3.4105
R787 VPWR.n164 VPWR.n163 3.4105
R788 VPWR.n236 VPWR.n235 3.4105
R789 VPWR.n674 VPWR.n673 3.4105
R790 VPWR.n674 VPWR.n54 3.4105
R791 VPWR.n673 VPWR.n672 3.4105
R792 VPWR.n62 VPWR.n54 3.4105
R793 VPWR.n129 VPWR.n128 3.4105
R794 VPWR.n130 VPWR.n56 3.4105
R795 VPWR.n527 VPWR.n525 3.4105
R796 VPWR.n585 VPWR.n584 3.4105
R797 VPWR.n75 VPWR.n74 3.4105
R798 VPWR.n99 VPWR.n98 3.4105
R799 VPWR.n207 VPWR.n206 3.4105
R800 VPWR.n206 VPWR.n205 3.4105
R801 VPWR.n208 VPWR.n207 3.4105
R802 VPWR.n205 VPWR.n204 3.4105
R803 VPWR.n180 VPWR.n178 3.4105
R804 VPWR.n199 VPWR.n176 3.4105
R805 VPWR.n622 VPWR.n621 3.4105
R806 VPWR.n599 VPWR.n280 3.4105
R807 VPWR.n431 VPWR.n430 3.4105
R808 VPWR.n431 VPWR.n282 3.4105
R809 VPWR.n430 VPWR.n429 3.4105
R810 VPWR.n408 VPWR.n282 3.4105
R811 VPWR.n411 VPWR.n410 3.4105
R812 VPWR.n412 VPWR.n283 3.4105
R813 VPWR.t49 VPWR.t199 3.35739
R814 VPWR.t144 VPWR.t31 3.35739
R815 VPWR.n25 VPWR.n24 3.05586
R816 VPWR.n85 VPWR.n84 3.05586
R817 VPWR.n190 VPWR.n189 3.05586
R818 VPWR.n506 VPWR.n505 3.04861
R819 VPWR.n580 VPWR.n579 3.04861
R820 VPWR.n613 VPWR.n612 3.04861
R821 VPWR.n455 VPWR.n451 3.01588
R822 VPWR.n489 VPWR.n488 3.01588
R823 VPWR.n659 VPWR.n142 3.01588
R824 VPWR.n557 VPWR.n556 3.01588
R825 VPWR.n42 VPWR.n39 2.8165
R826 VPWR.n458 VPWR.n451 2.64665
R827 VPWR.n490 VPWR.n489 2.64665
R828 VPWR.n538 VPWR.n142 2.64665
R829 VPWR.n20 VPWR.n18 2.63539
R830 VPWR.n23 VPWR.n21 2.63539
R831 VPWR.n501 VPWR.n499 2.63539
R832 VPWR.n504 VPWR.n502 2.63539
R833 VPWR.n80 VPWR.n78 2.63539
R834 VPWR.n83 VPWR.n81 2.63539
R835 VPWR.n575 VPWR.n573 2.63539
R836 VPWR.n578 VPWR.n576 2.63539
R837 VPWR.n185 VPWR.n183 2.63539
R838 VPWR.n188 VPWR.n186 2.63539
R839 VPWR.n608 VPWR.n606 2.63539
R840 VPWR.n611 VPWR.n609 2.63539
R841 VPWR.n22 VPWR.n21 2.37495
R842 VPWR.n19 VPWR.n18 2.37495
R843 VPWR.n503 VPWR.n502 2.37495
R844 VPWR.n500 VPWR.n499 2.37495
R845 VPWR.n82 VPWR.n81 2.37495
R846 VPWR.n79 VPWR.n78 2.37495
R847 VPWR.n577 VPWR.n576 2.37495
R848 VPWR.n574 VPWR.n573 2.37495
R849 VPWR.n187 VPWR.n186 2.37495
R850 VPWR.n184 VPWR.n183 2.37495
R851 VPWR.n610 VPWR.n609 2.37495
R852 VPWR.n607 VPWR.n606 2.37495
R853 VPWR.n371 VPWR.n370 2.33701
R854 VPWR.n696 VPWR.n694 2.29615
R855 VPWR.n556 VPWR.n532 2.27742
R856 VPWR.n705 VPWR.n704 2.25932
R857 VPWR.n632 VPWR.n273 2.25932
R858 VPWR.n370 VPWR.n369 2.03225
R859 VPWR.n668 VPWR.n667 1.85065
R860 VPWR.n138 VPWR.n137 1.69962
R861 VPWR.n653 VPWR.n148 1.69188
R862 VPWR.n653 VPWR.n652 1.69188
R863 VPWR.n654 VPWR.n147 1.69188
R864 VPWR.n655 VPWR.n654 1.69188
R865 VPWR.n390 VPWR.n389 1.69188
R866 VPWR.n389 VPWR.n388 1.69188
R867 VPWR.n474 VPWR.n146 1.69188
R868 VPWR.n237 VPWR.n55 1.69188
R869 VPWR.n225 VPWR.n55 1.69188
R870 VPWR.n683 VPWR.n682 1.69188
R871 VPWR.n682 VPWR.n681 1.69188
R872 VPWR.n358 VPWR.n52 1.69188
R873 VPWR.n355 VPWR.n52 1.69188
R874 VPWR.n674 VPWR.n53 1.69188
R875 VPWR.n100 VPWR.n8 1.69188
R876 VPWR.n88 VPWR.n8 1.69188
R877 VPWR.n718 VPWR.n7 1.69188
R878 VPWR.n718 VPWR.n717 1.69188
R879 VPWR.n719 VPWR.n6 1.69188
R880 VPWR.n720 VPWR.n719 1.69188
R881 VPWR.n206 VPWR.n177 1.69188
R882 VPWR.n619 VPWR.n618 1.69188
R883 VPWR.n620 VPWR.n619 1.69188
R884 VPWR.n598 VPWR.n524 1.69188
R885 VPWR.n598 VPWR.n597 1.69188
R886 VPWR.n523 VPWR.n432 1.69188
R887 VPWR.n523 VPWR.n522 1.69188
R888 VPWR.n431 VPWR.n281 1.69188
R889 VPWR.t35 VPWR.t107 1.67895
R890 VPWR.t121 VPWR.t37 1.67895
R891 VPWR.n137 VPWR.n136 1.54858
R892 VPWR.n667 VPWR.n666 1.39755
R893 VPWR.n694 VPWR.n693 1.36405
R894 VPWR.n216 VPWR.n215 1.12991
R895 VPWR.n43 VPWR.n42 1.11173
R896 VPWR.n420 VPWR.n418 0.863992
R897 VPWR.n322 VPWR.n2 0.863992
R898 VPWR.n727 VPWR.n726 0.863992
R899 VPWR.n565 VPWR.n564 0.833988
R900 VPWR.n254 VPWR.n253 0.833988
R901 VPWR.n32 VPWR.n31 0.753441
R902 VPWR.n93 VPWR.n92 0.635211
R903 VPWR.n106 VPWR.n105 0.635211
R904 VPWR.n581 VPWR.n571 0.635211
R905 VPWR.n231 VPWR.n160 0.635211
R906 VPWR.n245 VPWR.n244 0.635211
R907 VPWR.n646 VPWR.n645 0.635211
R908 VPWR.n378 VPWR.n377 0.635211
R909 VPWR.n404 VPWR.n403 0.635211
R910 VPWR.n568 VPWR.n530 0.595849
R911 VPWR.n250 VPWR.n154 0.595849
R912 VPWR.n688 VPWR.n46 0.369731
R913 VPWR.n481 VPWR.n442 0.369731
R914 VPWR.n483 VPWR.n482 0.369731
R915 VPWR.n507 VPWR.n497 0.369731
R916 VPWR.n141 VPWR.n139 0.369731
R917 VPWR.n550 VPWR.n536 0.369731
R918 VPWR.n551 VPWR.n534 0.369731
R919 VPWR.n560 VPWR.n532 0.369731
R920 VPWR.n630 VPWR.n274 0.305262
R921 VPWR.n614 VPWR.n605 0.305262
R922 VPWR.n425 VPWR.n418 0.305262
R923 VPWR.n369 VPWR.n368 0.305262
R924 VPWR.n372 VPWR.n304 0.305262
R925 VPWR.n724 VPWR.n2 0.305262
R926 VPWR.n325 VPWR.n324 0.305262
R927 VPWR.n726 VPWR.n725 0.305262
R928 VPWR.n26 VPWR.n25 0.232472
R929 VPWR.n86 VPWR.n85 0.232472
R930 VPWR.n191 VPWR.n190 0.232472
R931 VPWR.n136 VPWR.n135 0.227049
R932 VPWR.n666 VPWR.n665 0.227049
R933 VPWR.n505 VPWR 0.217591
R934 VPWR.n94 VPWR.n71 0.21207
R935 VPWR.n592 VPWR.n591 0.21207
R936 VPWR.n242 VPWR.n241 0.21207
R937 VPWR.n260 VPWR.n259 0.21207
R938 VPWR.n579 VPWR 0.208476
R939 VPWR.n612 VPWR 0.207174
R940 VPWR.n389 VPWR.n146 0.1603
R941 VPWR.n654 VPWR.n146 0.1603
R942 VPWR.n654 VPWR.n653 0.1603
R943 VPWR.n682 VPWR.n52 0.1603
R944 VPWR.n682 VPWR.n674 0.1603
R945 VPWR.n674 VPWR.n55 0.1603
R946 VPWR.n719 VPWR.n718 0.1603
R947 VPWR.n718 VPWR.n8 0.1603
R948 VPWR.n206 VPWR.n8 0.1603
R949 VPWR.n523 VPWR.n431 0.1603
R950 VPWR.n598 VPWR.n523 0.1603
R951 VPWR.n619 VPWR.n598 0.1603
R952 VPWR.n691 VPWR 0.159471
R953 VPWR VPWR.n698 0.149054
R954 VPWR.n505 VPWR 0.141725
R955 VPWR.n579 VPWR 0.141725
R956 VPWR.n612 VPWR 0.141725
R957 VPWR.n703 VPWR.n702 0.120292
R958 VPWR.n456 VPWR.n452 0.120292
R959 VPWR.n457 VPWR.n456 0.120292
R960 VPWR.n457 VPWR.n450 0.120292
R961 VPWR.n461 VPWR.n450 0.120292
R962 VPWR.n462 VPWR.n461 0.120292
R963 VPWR.n464 VPWR.n462 0.120292
R964 VPWR.n485 VPWR.n441 0.120292
R965 VPWR.n486 VPWR.n485 0.120292
R966 VPWR.n487 VPWR.n486 0.120292
R967 VPWR.n487 VPWR.n439 0.120292
R968 VPWR.n492 VPWR.n439 0.120292
R969 VPWR.n493 VPWR.n492 0.120292
R970 VPWR.n494 VPWR.n493 0.120292
R971 VPWR.n109 VPWR.n68 0.120292
R972 VPWR.n111 VPWR.n110 0.120292
R973 VPWR.n111 VPWR.n65 0.120292
R974 VPWR.n117 VPWR.n65 0.120292
R975 VPWR.n118 VPWR.n117 0.120292
R976 VPWR.n670 VPWR.n59 0.120292
R977 VPWR.n664 VPWR.n59 0.120292
R978 VPWR.n663 VPWR.n662 0.120292
R979 VPWR.n662 VPWR.n140 0.120292
R980 VPWR.n658 VPWR.n140 0.120292
R981 VPWR.n553 VPWR.n552 0.120292
R982 VPWR.n553 VPWR.n533 0.120292
R983 VPWR.n558 VPWR.n533 0.120292
R984 VPWR.n559 VPWR.n558 0.120292
R985 VPWR.n566 VPWR.n531 0.120292
R986 VPWR.n567 VPWR.n566 0.120292
R987 VPWR.n211 VPWR.n210 0.120292
R988 VPWR.n217 VPWR.n170 0.120292
R989 VPWR.n218 VPWR.n217 0.120292
R990 VPWR.n218 VPWR.n167 0.120292
R991 VPWR.n222 VPWR.n167 0.120292
R992 VPWR.n246 VPWR.n157 0.120292
R993 VPWR.n247 VPWR.n246 0.120292
R994 VPWR.n255 VPWR.n155 0.120292
R995 VPWR.n256 VPWR.n255 0.120292
R996 VPWR.n257 VPWR.n256 0.120292
R997 VPWR.n634 VPWR.n267 0.120292
R998 VPWR.n634 VPWR.n633 0.120292
R999 VPWR.n633 VPWR.n271 0.120292
R1000 VPWR.n629 VPWR.n628 0.120292
R1001 VPWR.n729 VPWR.n1 0.120292
R1002 VPWR.n723 VPWR.n1 0.120292
R1003 VPWR.n340 VPWR.n339 0.120292
R1004 VPWR.n341 VPWR.n340 0.120292
R1005 VPWR.n341 VPWR.n318 0.120292
R1006 VPWR.n345 VPWR.n318 0.120292
R1007 VPWR.n347 VPWR.n346 0.120292
R1008 VPWR.n366 VPWR.n365 0.120292
R1009 VPWR.n367 VPWR 0.120292
R1010 VPWR.n374 VPWR 0.120292
R1011 VPWR.n375 VPWR.n374 0.120292
R1012 VPWR.n394 VPWR.n393 0.120292
R1013 VPWR.n394 VPWR.n292 0.120292
R1014 VPWR.n398 VPWR.n292 0.120292
R1015 VPWR.n399 VPWR.n398 0.120292
R1016 VPWR.n400 VPWR.n399 0.120292
R1017 VPWR.n400 VPWR.n290 0.120292
R1018 VPWR.n405 VPWR.n290 0.120292
R1019 VPWR.n424 VPWR.n423 0.120292
R1020 VPWR.n423 VPWR.n419 0.120292
R1021 VPWR.n464 VPWR.n463 0.11899
R1022 VPWR.n658 VPWR.n657 0.11899
R1023 VPWR.n257 VPWR.n150 0.11899
R1024 VPWR.n376 VPWR.n298 0.11899
R1025 VPWR.n452 VPWR.n50 0.117688
R1026 VPWR.n671 VPWR.n670 0.117688
R1027 VPWR.n239 VPWR.n157 0.117688
R1028 VPWR.n365 VPWR.n306 0.117688
R1029 VPWR.n25 VPWR 0.105238
R1030 VPWR.n85 VPWR 0.105238
R1031 VPWR.n190 VPWR 0.105238
R1032 VPWR.n346 VPWR 0.0994583
R1033 VPWR.n699 VPWR 0.0981562
R1034 VPWR VPWR.n690 0.0981562
R1035 VPWR.n110 VPWR 0.0981562
R1036 VPWR.n120 VPWR 0.0981562
R1037 VPWR VPWR.n663 0.0981562
R1038 VPWR VPWR.n531 0.0981562
R1039 VPWR VPWR.n170 0.0981562
R1040 VPWR.n223 VPWR 0.0981562
R1041 VPWR VPWR.n155 0.0981562
R1042 VPWR.n629 VPWR 0.0981562
R1043 VPWR VPWR.n729 0.0981562
R1044 VPWR.n376 VPWR 0.0981562
R1045 VPWR.n424 VPWR 0.0981562
R1046 VPWR.n267 VPWR 0.0968542
R1047 VPWR.n721 VPWR.n4 0.0950946
R1048 VPWR.n334 VPWR.n333 0.0950946
R1049 VPWR.n354 VPWR.n353 0.0950946
R1050 VPWR.n360 VPWR.n359 0.0950946
R1051 VPWR.n387 VPWR.n386 0.0950946
R1052 VPWR.n391 VPWR.n295 0.0950946
R1053 VPWR.n656 VPWR.n144 0.0950946
R1054 VPWR.n547 VPWR.n546 0.0950946
R1055 VPWR.n651 VPWR.n650 0.0950946
R1056 VPWR.n642 VPWR.n641 0.0950946
R1057 VPWR.n470 VPWR.n447 0.0950946
R1058 VPWR.n478 VPWR.n477 0.0950946
R1059 VPWR.n716 VPWR.n715 0.0950946
R1060 VPWR.n709 VPWR.n14 0.0950946
R1061 VPWR.n521 VPWR.n520 0.0950946
R1062 VPWR.n513 VPWR.n512 0.0950946
R1063 VPWR.n680 VPWR.n679 0.0950946
R1064 VPWR.n685 VPWR.n684 0.0950946
R1065 VPWR.n227 VPWR.n226 0.0950946
R1066 VPWR.n238 VPWR.n162 0.0950946
R1067 VPWR.n127 VPWR.n62 0.0950946
R1068 VPWR.n672 VPWR.n57 0.0950946
R1069 VPWR.n596 VPWR.n595 0.0950946
R1070 VPWR.n587 VPWR.n586 0.0950946
R1071 VPWR.n89 VPWR.n87 0.0950946
R1072 VPWR.n101 VPWR.n73 0.0950946
R1073 VPWR.n204 VPWR.n203 0.0950946
R1074 VPWR.n208 VPWR.n175 0.0950946
R1075 VPWR.n623 VPWR.n278 0.0950946
R1076 VPWR.n617 VPWR.n600 0.0950946
R1077 VPWR.n409 VPWR.n408 0.0950946
R1078 VPWR.n429 VPWR.n284 0.0950946
R1079 VPWR.n494 VPWR.n434 0.0890417
R1080 VPWR.n567 VPWR.n526 0.0890417
R1081 VPWR.n628 VPWR.n275 0.0890417
R1082 VPWR.n367 VPWR 0.0890417
R1083 VPWR.n703 VPWR.n15 0.0877396
R1084 VPWR.n102 VPWR.n68 0.0877396
R1085 VPWR.n210 VPWR.n209 0.0877396
R1086 VPWR VPWR.n638 0.0877396
R1087 VPWR.n339 VPWR.n320 0.0877396
R1088 VPWR VPWR.n315 0.0877396
R1089 VPWR.n653 VPWR 0.08745
R1090 VPWR.n55 VPWR 0.08745
R1091 VPWR.n206 VPWR 0.08745
R1092 VPWR.n619 VPWR 0.08745
R1093 VPWR.n714 VPWR.n713 0.0838333
R1094 VPWR.n498 VPWR.n437 0.0838333
R1095 VPWR.n96 VPWR.n76 0.0838333
R1096 VPWR.n572 VPWR.n529 0.0838333
R1097 VPWR.n202 VPWR.n201 0.0838333
R1098 VPWR.n602 VPWR.n601 0.0838333
R1099 VPWR.n329 VPWR.n327 0.0838333
R1100 VPWR.n392 VPWR.n294 0.0838333
R1101 VPWR.n414 VPWR.n289 0.0838333
R1102 VPWR.n691 VPWR 0.082648
R1103 VPWR.n469 VPWR.n448 0.0825312
R1104 VPWR.n537 VPWR.n143 0.0825312
R1105 VPWR.n649 VPWR.n152 0.0825312
R1106 VPWR.n385 VPWR.n300 0.0825312
R1107 VPWR.n698 VPWR 0.0813459
R1108 VPWR.n678 VPWR 0.0812292
R1109 VPWR.n686 VPWR.n48 0.0812292
R1110 VPWR.n126 VPWR 0.0812292
R1111 VPWR.n133 VPWR.n58 0.0812292
R1112 VPWR.n228 VPWR 0.0812292
R1113 VPWR.n240 VPWR.n161 0.0812292
R1114 VPWR.n352 VPWR 0.0812292
R1115 VPWR.n362 VPWR.n361 0.0812292
R1116 VPWR.n480 VPWR.n443 0.0747188
R1117 VPWR.n549 VPWR.n541 0.0747188
R1118 VPWR.n644 VPWR.n262 0.0747188
R1119 VPWR.n381 VPWR.n303 0.0747188
R1120 VPWR.n445 VPWR 0.0708125
R1121 VPWR VPWR.n535 0.0708125
R1122 VPWR.n640 VPWR 0.0708125
R1123 VPWR.n708 VPWR.n13 0.0695104
R1124 VPWR.n95 VPWR.n72 0.0695104
R1125 VPWR.n198 VPWR.n182 0.0695104
R1126 VPWR.n519 VPWR.n518 0.0682083
R1127 VPWR.n594 VPWR.n593 0.0682083
R1128 VPWR.n624 VPWR.n277 0.0682083
R1129 VPWR.n415 VPWR.n288 0.0682083
R1130 VPWR.n330 VPWR.n326 0.0680676
R1131 VPWR.n332 VPWR.n330 0.0680676
R1132 VPWR.n313 VPWR.n311 0.0680676
R1133 VPWR.n313 VPWR.n310 0.0680676
R1134 VPWR.n302 VPWR.n299 0.0680676
R1135 VPWR.n302 VPWR.n301 0.0680676
R1136 VPWR.n543 VPWR.n542 0.0680676
R1137 VPWR.n545 VPWR.n543 0.0680676
R1138 VPWR.n263 VPWR.n151 0.0680676
R1139 VPWR.n265 VPWR.n263 0.0680676
R1140 VPWR.n472 VPWR.n471 0.0680676
R1141 VPWR.n471 VPWR.n444 0.0680676
R1142 VPWR.n712 VPWR.n11 0.0680676
R1143 VPWR.n712 VPWR.n711 0.0680676
R1144 VPWR.n509 VPWR.n435 0.0680676
R1145 VPWR.n511 VPWR.n509 0.0680676
R1146 VPWR.n677 VPWR.n676 0.0680676
R1147 VPWR.n676 VPWR.n49 0.0680676
R1148 VPWR.n234 VPWR.n164 0.0680676
R1149 VPWR.n235 VPWR.n234 0.0680676
R1150 VPWR.n131 VPWR.n129 0.0680676
R1151 VPWR.n131 VPWR.n130 0.0680676
R1152 VPWR.n583 VPWR.n527 0.0680676
R1153 VPWR.n585 VPWR.n583 0.0680676
R1154 VPWR.n97 VPWR.n75 0.0680676
R1155 VPWR.n98 VPWR.n97 0.0680676
R1156 VPWR.n200 VPWR.n180 0.0680676
R1157 VPWR.n200 VPWR.n199 0.0680676
R1158 VPWR.n622 VPWR.n279 0.0680676
R1159 VPWR.n599 VPWR.n279 0.0680676
R1160 VPWR.n413 VPWR.n411 0.0680676
R1161 VPWR.n413 VPWR.n412 0.0680676
R1162 VPWR.n407 VPWR 0.0669062
R1163 VPWR.n515 VPWR.n514 0.063
R1164 VPWR.n616 VPWR.n603 0.063
R1165 VPWR.n428 VPWR.n285 0.063
R1166 VPWR.n12 VPWR.n10 0.0616979
R1167 VPWR.n91 VPWR.n90 0.0616979
R1168 VPWR.n181 VPWR.n179 0.0616979
R1169 VPWR.n722 VPWR.n3 0.0616979
R1170 VPWR.n26 VPWR.n10 0.0590938
R1171 VPWR.n191 VPWR.n179 0.0590938
R1172 VPWR.n723 VPWR.n722 0.0590938
R1173 VPWR.n514 VPWR.n508 0.0577917
R1174 VPWR.n588 VPWR.n582 0.0577917
R1175 VPWR.n616 VPWR.n615 0.0577917
R1176 VPWR.n428 VPWR.n427 0.0577917
R1177 VPWR.n331 VPWR.n5 0.0574697
R1178 VPWR.n357 VPWR.n356 0.0574697
R1179 VPWR.n297 VPWR.n296 0.0574697
R1180 VPWR.n544 VPWR.n145 0.0574697
R1181 VPWR.n264 VPWR.n149 0.0574697
R1182 VPWR.n473 VPWR.n446 0.0574697
R1183 VPWR.n476 VPWR.n475 0.0574697
R1184 VPWR.n710 VPWR.n9 0.0574697
R1185 VPWR.n510 VPWR.n433 0.0574697
R1186 VPWR.n675 VPWR.n51 0.0574697
R1187 VPWR.n236 VPWR.n163 0.0574697
R1188 VPWR.n128 VPWR.n54 0.0574697
R1189 VPWR.n673 VPWR.n56 0.0574697
R1190 VPWR.n584 VPWR.n525 0.0574697
R1191 VPWR.n99 VPWR.n74 0.0574697
R1192 VPWR.n205 VPWR.n178 0.0574697
R1193 VPWR.n207 VPWR.n176 0.0574697
R1194 VPWR.n621 VPWR.n280 0.0574697
R1195 VPWR.n410 VPWR.n282 0.0574697
R1196 VPWR.n430 VPWR.n283 0.0574697
R1197 VPWR.n132 VPWR 0.0538854
R1198 VPWR VPWR.n314 0.0538854
R1199 VPWR.n519 VPWR.n436 0.0525833
R1200 VPWR.n594 VPWR.n528 0.0525833
R1201 VPWR.n625 VPWR.n624 0.0525833
R1202 VPWR.n406 VPWR.n288 0.0525833
R1203 VPWR.n708 VPWR.n707 0.0512812
R1204 VPWR.n103 VPWR.n72 0.0512812
R1205 VPWR.n182 VPWR.n174 0.0512812
R1206 VPWR.n336 VPWR.n335 0.0512812
R1207 VPWR.n335 VPWR 0.047375
R1208 VPWR.n468 VPWR.n443 0.0460729
R1209 VPWR.n541 VPWR.n540 0.0460729
R1210 VPWR.n384 VPWR.n303 0.0460729
R1211 VPWR.n47 VPWR 0.0447708
R1212 VPWR.n687 VPWR.n47 0.0447708
R1213 VPWR.n134 VPWR.n132 0.0447708
R1214 VPWR.n233 VPWR 0.0447708
R1215 VPWR.n233 VPWR.n232 0.0447708
R1216 VPWR.n314 VPWR.n309 0.0447708
R1217 VPWR.n326 VPWR.n4 0.0410405
R1218 VPWR.n334 VPWR.n332 0.0410405
R1219 VPWR.n353 VPWR.n311 0.0410405
R1220 VPWR.n360 VPWR.n310 0.0410405
R1221 VPWR.n386 VPWR.n299 0.0410405
R1222 VPWR.n301 VPWR.n295 0.0410405
R1223 VPWR.n542 VPWR.n144 0.0410405
R1224 VPWR.n547 VPWR.n545 0.0410405
R1225 VPWR.n650 VPWR.n151 0.0410405
R1226 VPWR.n642 VPWR.n265 0.0410405
R1227 VPWR.n472 VPWR.n470 0.0410405
R1228 VPWR.n478 VPWR.n444 0.0410405
R1229 VPWR.n715 VPWR.n11 0.0410405
R1230 VPWR.n711 VPWR.n709 0.0410405
R1231 VPWR.n520 VPWR.n435 0.0410405
R1232 VPWR.n512 VPWR.n511 0.0410405
R1233 VPWR.n679 VPWR.n677 0.0410405
R1234 VPWR.n685 VPWR.n49 0.0410405
R1235 VPWR.n227 VPWR.n164 0.0410405
R1236 VPWR.n235 VPWR.n162 0.0410405
R1237 VPWR.n129 VPWR.n127 0.0410405
R1238 VPWR.n130 VPWR.n57 0.0410405
R1239 VPWR.n595 VPWR.n527 0.0410405
R1240 VPWR.n586 VPWR.n585 0.0410405
R1241 VPWR.n87 VPWR.n75 0.0410405
R1242 VPWR.n98 VPWR.n73 0.0410405
R1243 VPWR.n203 VPWR.n180 0.0410405
R1244 VPWR.n199 VPWR.n175 0.0410405
R1245 VPWR.n623 VPWR.n622 0.0410405
R1246 VPWR.n600 VPWR.n599 0.0410405
R1247 VPWR.n411 VPWR.n409 0.0410405
R1248 VPWR.n412 VPWR.n284 0.0410405
R1249 VPWR VPWR.n588 0.0408646
R1250 VPWR.n687 VPWR.n686 0.0395625
R1251 VPWR.n134 VPWR.n133 0.0395625
R1252 VPWR.n232 VPWR.n161 0.0395625
R1253 VPWR.n361 VPWR.n309 0.0395625
R1254 VPWR.n469 VPWR.n468 0.0382604
R1255 VPWR.n540 VPWR.n537 0.0382604
R1256 VPWR.n649 VPWR.n648 0.0382604
R1257 VPWR.n385 VPWR.n384 0.0382604
R1258 VPWR.n707 VPWR.n15 0.0330521
R1259 VPWR.n103 VPWR.n102 0.0330521
R1260 VPWR.n209 VPWR.n174 0.0330521
R1261 VPWR.n639 VPWR 0.0330521
R1262 VPWR.n336 VPWR.n320 0.0330521
R1263 VPWR.n347 VPWR 0.0330521
R1264 VPWR.n699 VPWR 0.03175
R1265 VPWR.n436 VPWR.n434 0.03175
R1266 VPWR VPWR.n86 0.03175
R1267 VPWR.n528 VPWR.n526 0.03175
R1268 VPWR.n229 VPWR 0.03175
R1269 VPWR.n625 VPWR.n275 0.03175
R1270 VPWR VPWR.n366 0.03175
R1271 VPWR.n407 VPWR.n406 0.03175
R1272 VPWR.n652 VPWR.n149 0.0292489
R1273 VPWR.n264 VPWR.n148 0.0292489
R1274 VPWR.n655 VPWR.n145 0.0292489
R1275 VPWR.n544 VPWR.n147 0.0292489
R1276 VPWR.n388 VPWR.n297 0.0292489
R1277 VPWR.n390 VPWR.n296 0.0292489
R1278 VPWR.n475 VPWR.n474 0.0292489
R1279 VPWR.n474 VPWR.n473 0.0292489
R1280 VPWR.n225 VPWR.n163 0.0292489
R1281 VPWR.n237 VPWR.n236 0.0292489
R1282 VPWR.n681 VPWR.n675 0.0292489
R1283 VPWR.n683 VPWR.n51 0.0292489
R1284 VPWR.n356 VPWR.n355 0.0292489
R1285 VPWR.n358 VPWR.n357 0.0292489
R1286 VPWR.n56 VPWR.n53 0.0292489
R1287 VPWR.n128 VPWR.n53 0.0292489
R1288 VPWR.n88 VPWR.n74 0.0292489
R1289 VPWR.n100 VPWR.n99 0.0292489
R1290 VPWR.n717 VPWR.n9 0.0292489
R1291 VPWR.n710 VPWR.n7 0.0292489
R1292 VPWR.n720 VPWR.n5 0.0292489
R1293 VPWR.n331 VPWR.n6 0.0292489
R1294 VPWR.n177 VPWR.n176 0.0292489
R1295 VPWR.n178 VPWR.n177 0.0292489
R1296 VPWR.n621 VPWR.n620 0.0292489
R1297 VPWR.n618 VPWR.n280 0.0292489
R1298 VPWR.n597 VPWR.n525 0.0292489
R1299 VPWR.n584 VPWR.n524 0.0292489
R1300 VPWR.n522 VPWR.n433 0.0292489
R1301 VPWR.n510 VPWR.n432 0.0292489
R1302 VPWR.n283 VPWR.n281 0.0292489
R1303 VPWR.n410 VPWR.n281 0.0292489
R1304 VPWR.n690 VPWR.n40 0.0291458
R1305 VPWR.n120 VPWR.n119 0.0291458
R1306 VPWR.n315 VPWR.n312 0.0291458
R1307 VPWR.n445 VPWR.n441 0.0278438
R1308 VPWR.n90 VPWR 0.0278438
R1309 VPWR.n552 VPWR.n535 0.0278438
R1310 VPWR.n640 VPWR.n639 0.0278438
R1311 VPWR.n393 VPWR.n392 0.0278438
R1312 VPWR.n262 VPWR 0.0239375
R1313 VPWR.n638 VPWR 0.0239375
R1314 VPWR.n714 VPWR.n12 0.0226354
R1315 VPWR.n702 VPWR 0.0226354
R1316 VPWR VPWR.n44 0.0226354
R1317 VPWR.n508 VPWR 0.0226354
R1318 VPWR.n91 VPWR.n76 0.0226354
R1319 VPWR VPWR.n109 0.0226354
R1320 VPWR VPWR.n118 0.0226354
R1321 VPWR.n125 VPWR 0.0226354
R1322 VPWR.n664 VPWR 0.0226354
R1323 VPWR.n559 VPWR 0.0226354
R1324 VPWR.n589 VPWR 0.0226354
R1325 VPWR.n582 VPWR 0.0226354
R1326 VPWR.n202 VPWR.n181 0.0226354
R1327 VPWR.n211 VPWR 0.0226354
R1328 VPWR VPWR.n222 0.0226354
R1329 VPWR.n247 VPWR 0.0226354
R1330 VPWR.n648 VPWR 0.0226354
R1331 VPWR VPWR.n271 0.0226354
R1332 VPWR.n615 VPWR 0.0226354
R1333 VPWR.n327 VPWR.n3 0.0226354
R1334 VPWR.n328 VPWR 0.0226354
R1335 VPWR.n351 VPWR 0.0226354
R1336 VPWR VPWR.n375 0.0226354
R1337 VPWR VPWR.n405 0.0226354
R1338 VPWR.n427 VPWR 0.0226354
R1339 VPWR.n419 VPWR 0.0226354
R1340 VPWR.n515 VPWR.n498 0.0213333
R1341 VPWR.n589 VPWR.n572 0.0213333
R1342 VPWR VPWR.n223 0.0213333
R1343 VPWR.n603 VPWR.n602 0.0213333
R1344 VPWR VPWR.n345 0.0213333
R1345 VPWR.n289 VPWR.n285 0.0213333
R1346 VPWR.n518 VPWR.n437 0.016125
R1347 VPWR.n593 VPWR.n529 0.016125
R1348 VPWR.n601 VPWR.n277 0.016125
R1349 VPWR.n415 VPWR.n414 0.016125
R1350 VPWR.n713 VPWR.n13 0.0148229
R1351 VPWR.n96 VPWR.n95 0.0148229
R1352 VPWR.n201 VPWR.n198 0.0148229
R1353 VPWR.n329 VPWR.n328 0.0148229
R1354 VPWR.n479 VPWR 0.0135208
R1355 VPWR.n548 VPWR 0.0135208
R1356 VPWR.n643 VPWR 0.0135208
R1357 VPWR.n480 VPWR.n479 0.00961458
R1358 VPWR.n549 VPWR.n548 0.00961458
R1359 VPWR.n644 VPWR.n643 0.00961458
R1360 VPWR.n381 VPWR.n294 0.00961458
R1361 VPWR.n678 VPWR.n44 0.0083125
R1362 VPWR.n126 VPWR.n125 0.0083125
R1363 VPWR.n224 VPWR 0.0083125
R1364 VPWR.n229 VPWR.n228 0.0083125
R1365 VPWR.n352 VPWR.n351 0.0083125
R1366 VPWR VPWR.n40 0.00310417
R1367 VPWR.n50 VPWR.n48 0.00310417
R1368 VPWR.n119 VPWR 0.00310417
R1369 VPWR.n671 VPWR.n58 0.00310417
R1370 VPWR.n224 VPWR 0.00310417
R1371 VPWR.n240 VPWR.n239 0.00310417
R1372 VPWR VPWR.n312 0.00310417
R1373 VPWR.n362 VPWR.n306 0.00310417
R1374 VPWR.n463 VPWR.n448 0.00180208
R1375 VPWR.n657 VPWR.n143 0.00180208
R1376 VPWR.n152 VPWR.n150 0.00180208
R1377 VPWR.n300 VPWR.n298 0.00180208
R1378 VGND.n305 VGND.n140 16191.9
R1379 VGND.n388 VGND 9498.47
R1380 VGND.n389 VGND.n140 4986.67
R1381 VGND.n389 VGND.n388 4986.67
R1382 VGND VGND.t165 4897.32
R1383 VGND VGND.t171 4888.89
R1384 VGND.t171 VGND 4408.43
R1385 VGND.t165 VGND 4408.43
R1386 VGND VGND.n307 3807.53
R1387 VGND.t126 VGND.t138 3101.92
R1388 VGND.n306 VGND.n305 2415.34
R1389 VGND.n307 VGND.n306 2415.34
R1390 VGND.t141 VGND.t174 2326.44
R1391 VGND.t121 VGND.t29 2022.99
R1392 VGND VGND.t126 1795.4
R1393 VGND VGND.t132 1786.97
R1394 VGND.t168 VGND 1702.68
R1395 VGND.t62 VGND.t1 1584.67
R1396 VGND.t199 VGND.t191 1550.96
R1397 VGND VGND.t160 1407.66
R1398 VGND VGND.t129 1407.66
R1399 VGND.t194 VGND 1399.23
R1400 VGND.t84 VGND 1340.23
R1401 VGND.t191 VGND 1306.51
R1402 VGND.t132 VGND 1306.51
R1403 VGND.t138 VGND 1306.51
R1404 VGND VGND.t150 1289.66
R1405 VGND.n387 VGND.n386 1198.25
R1406 VGND.n644 VGND.n78 1198.25
R1407 VGND.n414 VGND.n390 1194.5
R1408 VGND.n304 VGND.n303 1194.5
R1409 VGND.t96 VGND.t90 1180.08
R1410 VGND.t33 VGND 1112.64
R1411 VGND VGND.t41 1053.64
R1412 VGND.t155 VGND 1047.19
R1413 VGND VGND.t80 1045.21
R1414 VGND.t14 VGND 1036.78
R1415 VGND VGND.t155 944.277
R1416 VGND.n390 VGND 918.774
R1417 VGND.t160 VGND 918.774
R1418 VGND VGND.t194 918.774
R1419 VGND.n304 VGND 918.774
R1420 VGND.t129 VGND 918.774
R1421 VGND.n306 VGND 851.341
R1422 VGND.n307 VGND 851.341
R1423 VGND.t59 VGND 851.341
R1424 VGND.n305 VGND 851.341
R1425 VGND.t107 VGND.t14 826.054
R1426 VGND.t12 VGND.t119 817.625
R1427 VGND.t27 VGND.t2 817.625
R1428 VGND.t202 VGND.t39 817.625
R1429 VGND.t4 VGND.t86 800.766
R1430 VGND.t82 VGND.t43 800.766
R1431 VGND.t6 VGND.t8 724.904
R1432 VGND.t8 VGND.t10 724.904
R1433 VGND.t10 VGND.t12 724.904
R1434 VGND.t29 VGND.t31 724.904
R1435 VGND.t31 VGND.t25 724.904
R1436 VGND.t25 VGND.t27 724.904
R1437 VGND.t35 VGND.t33 724.904
R1438 VGND.t37 VGND.t35 724.904
R1439 VGND.t39 VGND.t182 708.047
R1440 VGND.t66 VGND.t52 708.047
R1441 VGND.t50 VGND.t66 708.047
R1442 VGND.t104 VGND.t46 708.047
R1443 VGND.t65 VGND.t56 708.047
R1444 VGND.t100 VGND.t113 708.047
R1445 VGND.t113 VGND.t94 708.047
R1446 VGND.t86 VGND.t84 708.047
R1447 VGND.t80 VGND.t82 708.047
R1448 VGND.t1 VGND.t107 657.471
R1449 VGND VGND.t168 632.184
R1450 VGND.n390 VGND 632.184
R1451 VGND VGND.t121 632.184
R1452 VGND VGND.t141 632.184
R1453 VGND VGND.t50 615.327
R1454 VGND.t45 VGND.t54 606.898
R1455 VGND.t88 VGND.t74 606.898
R1456 VGND VGND.n389 564.751
R1457 VGND.n388 VGND 564.751
R1458 VGND VGND.t64 564.751
R1459 VGND VGND.n140 564.751
R1460 VGND.t119 VGND 556.322
R1461 VGND.t2 VGND 556.322
R1462 VGND VGND.t202 556.322
R1463 VGND.t144 VGND 550.678
R1464 VGND VGND.t62 547.894
R1465 VGND VGND.t96 547.894
R1466 VGND.t43 VGND 547.894
R1467 VGND.t94 VGND 539.465
R1468 VGND.t64 VGND.t72 488.889
R1469 VGND.t68 VGND.t111 472.031
R1470 VGND.t92 VGND.t204 472.031
R1471 VGND VGND.t144 445.959
R1472 VGND.t111 VGND.t109 438.315
R1473 VGND.t206 VGND.t59 438.315
R1474 VGND.t212 VGND.t147 433.32
R1475 VGND.t57 VGND.n78 404.599
R1476 VGND.t90 VGND.t0 404.599
R1477 VGND.t179 VGND.n304 387.74
R1478 VGND.t41 VGND.t68 354.024
R1479 VGND.t48 VGND.t92 354.024
R1480 VGND.t102 VGND.t48 354.024
R1481 VGND.t70 VGND 334.017
R1482 VGND VGND.t6 320.307
R1483 VGND.t0 VGND.t102 303.449
R1484 VGND.t135 VGND 301.519
R1485 VGND.t52 VGND 286.591
R1486 VGND.n542 VGND.t91 280.978
R1487 VGND.n282 VGND.t234 276.115
R1488 VGND.t109 VGND.t206 269.733
R1489 VGND.n254 VGND.t237 265.298
R1490 VGND.n11 VGND.t226 262.784
R1491 VGND.n19 VGND.t228 262.784
R1492 VGND.n470 VGND.t231 262.784
R1493 VGND.n471 VGND.t233 262.784
R1494 VGND.n45 VGND.t217 262.784
R1495 VGND.n46 VGND.t219 262.784
R1496 VGND.n533 VGND.t220 262.784
R1497 VGND.n534 VGND.t222 262.784
R1498 VGND.n157 VGND.t235 262.784
R1499 VGND.n159 VGND.t236 262.784
R1500 VGND.n242 VGND.t240 262.784
R1501 VGND.n244 VGND.t242 262.784
R1502 VGND.n408 VGND.t245 262.719
R1503 VGND.n129 VGND.t225 262.719
R1504 VGND.n129 VGND.t224 262.719
R1505 VGND.n481 VGND.t230 262.719
R1506 VGND.n481 VGND.t227 262.719
R1507 VGND.n109 VGND.t238 262.719
R1508 VGND.n516 VGND.t239 262.719
R1509 VGND.n225 VGND.t218 262.719
R1510 VGND VGND.t179 261.303
R1511 VGND VGND.t4 261.303
R1512 VGND.n338 VGND.t241 259.082
R1513 VGND.n582 VGND.t244 259.082
R1514 VGND.n163 VGND.t232 259.082
R1515 VGND.n370 VGND.t99 246.506
R1516 VGND.t150 VGND 244.445
R1517 VGND.n681 VGND.t7 243.286
R1518 VGND.n320 VGND.t213 243.286
R1519 VGND.n604 VGND.t24 243.286
R1520 VGND.n43 VGND.t115 243.286
R1521 VGND.n43 VGND.t30 243.286
R1522 VGND.n532 VGND.t97 240.575
R1523 VGND.n81 VGND.t34 239.4
R1524 VGND.n501 VGND.t63 237.327
R1525 VGND.t23 VGND 236.52
R1526 VGND VGND.t199 236.016
R1527 VGND.t204 VGND.t104 236.016
R1528 VGND VGND.t57 227.587
R1529 VGND.t72 VGND.t45 219.157
R1530 VGND.n409 VGND.t223 218.308
R1531 VGND.n142 VGND.t221 218.308
R1532 VGND.n218 VGND.t216 218.308
R1533 VGND.n475 VGND.t186 214.456
R1534 VGND.n451 VGND.t185 214.456
R1535 VGND.n475 VGND.t167 214.456
R1536 VGND.n451 VGND.t166 214.456
R1537 VGND.n445 VGND.t190 214.456
R1538 VGND.n419 VGND.t189 214.456
R1539 VGND.n445 VGND.t173 214.456
R1540 VGND.n419 VGND.t172 214.456
R1541 VGND.n139 VGND.t201 214.456
R1542 VGND.n391 VGND.t193 214.456
R1543 VGND.n393 VGND.t192 214.456
R1544 VGND.n20 VGND.t200 214.456
R1545 VGND.n11 VGND.t188 214.456
R1546 VGND.n11 VGND.t187 214.456
R1547 VGND.n19 VGND.t170 214.456
R1548 VGND.n19 VGND.t169 214.456
R1549 VGND.n470 VGND.t178 214.456
R1550 VGND.n470 VGND.t177 214.456
R1551 VGND.n471 VGND.t162 214.456
R1552 VGND.n471 VGND.t161 214.456
R1553 VGND.n581 VGND.t137 214.456
R1554 VGND.n584 VGND.t136 214.456
R1555 VGND.n576 VGND.t146 214.456
R1556 VGND.n591 VGND.t145 214.456
R1557 VGND.n110 VGND.t157 214.456
R1558 VGND.n377 VGND.t156 214.456
R1559 VGND.n340 VGND.t149 214.456
R1560 VGND.n337 VGND.t148 214.456
R1561 VGND.n45 VGND.t123 214.456
R1562 VGND.n45 VGND.t122 214.456
R1563 VGND.n46 VGND.t125 214.456
R1564 VGND.n46 VGND.t124 214.456
R1565 VGND.n524 VGND.t152 214.456
R1566 VGND.n87 VGND.t151 214.456
R1567 VGND.n83 VGND.t184 214.456
R1568 VGND.n80 VGND.t183 214.456
R1569 VGND.n533 VGND.t196 214.456
R1570 VGND.n533 VGND.t195 214.456
R1571 VGND.n534 VGND.t198 214.456
R1572 VGND.n534 VGND.t197 214.456
R1573 VGND.n256 VGND.t128 214.456
R1574 VGND.n224 VGND.t139 214.456
R1575 VGND.n220 VGND.t127 214.456
R1576 VGND.n276 VGND.t154 214.456
R1577 VGND.n219 VGND.t134 214.456
R1578 VGND.n207 VGND.t133 214.456
R1579 VGND.n197 VGND.t153 214.456
R1580 VGND.n196 VGND.t181 214.456
R1581 VGND.n192 VGND.t180 214.456
R1582 VGND.n155 VGND.t176 214.456
R1583 VGND.n162 VGND.t175 214.456
R1584 VGND.n157 VGND.t164 214.456
R1585 VGND.n157 VGND.t163 214.456
R1586 VGND.n159 VGND.t143 214.456
R1587 VGND.n159 VGND.t142 214.456
R1588 VGND.n247 VGND.t140 214.456
R1589 VGND.n242 VGND.t159 214.456
R1590 VGND.n242 VGND.t158 214.456
R1591 VGND.n244 VGND.t131 214.456
R1592 VGND.n244 VGND.t130 214.456
R1593 VGND.n311 VGND.n310 210.601
R1594 VGND.n522 VGND.n498 207.965
R1595 VGND.n526 VGND.n497 207.965
R1596 VGND.n531 VGND.n530 207.965
R1597 VGND.n145 VGND.n144 207.213
R1598 VGND.n173 VGND.n152 207.213
R1599 VGND.n347 VGND.n346 205.078
R1600 VGND.n113 VGND.n112 205.078
R1601 VGND.n65 VGND.n41 205.078
R1602 VGND.n65 VGND.n42 205.078
R1603 VGND.n318 VGND.n317 203.619
R1604 VGND.n574 VGND.n566 203.619
R1605 VGND.n39 VGND.n37 203.619
R1606 VGND.n39 VGND.n38 203.619
R1607 VGND.n676 VGND.n22 200.812
R1608 VGND.n638 VGND.n82 200.812
R1609 VGND.n636 VGND.n86 200.561
R1610 VGND.n659 VGND.n73 200.105
R1611 VGND.n674 VGND.n23 199.662
R1612 VGND VGND.n387 198.606
R1613 VGND.n154 VGND.n153 198.475
R1614 VGND.n504 VGND.n503 197.476
R1615 VGND.n528 VGND.n527 197.476
R1616 VGND VGND.t135 196.799
R1617 VGND.n200 VGND.n199 196.442
R1618 VGND.n241 VGND.n240 196.442
R1619 VGND.n660 VGND.n72 195.612
R1620 VGND.n647 VGND.n646 185
R1621 VGND.n645 VGND.n74 185
R1622 VGND.n174 VGND.n145 185
R1623 VGND.n176 VGND.n175 185
R1624 VGND.t78 VGND.t210 175.133
R1625 VGND.t60 VGND.t70 175.133
R1626 VGND.t76 VGND.t21 175.133
R1627 VGND VGND.t98 169.718
R1628 VGND.t214 VGND.t212 155.274
R1629 VGND.t208 VGND.t214 155.274
R1630 VGND.t210 VGND.t208 155.274
R1631 VGND.t17 VGND.t23 155.274
R1632 VGND.t19 VGND.t17 155.274
R1633 VGND.t21 VGND.t19 155.274
R1634 VGND.t98 VGND.t60 151.662
R1635 VGND.n294 VGND.t85 150.376
R1636 VGND.n253 VGND.t81 150.376
R1637 VGND.n499 VGND.t53 146.964
R1638 VGND.t56 VGND 143.296
R1639 VGND.n646 VGND.n645 137.143
R1640 VGND.n175 VGND.n174 137.143
R1641 VGND.t147 VGND 135.412
R1642 VGND.n387 VGND 135.412
R1643 VGND VGND.n78 134.867
R1644 VGND.n576 VGND.t243 121.927
R1645 VGND.n83 VGND.t229 121.927
R1646 VGND VGND.t78 119.163
R1647 VGND VGND.t76 119.163
R1648 VGND.t54 VGND.t88 101.15
R1649 VGND.t74 VGND.t100 101.15
R1650 VGND.t46 VGND 92.7208
R1651 VGND.n73 VGND.t110 72.8576
R1652 VGND.t174 VGND.t65 67.4335
R1653 VGND.n503 VGND.t108 58.5719
R1654 VGND.n527 VGND.t49 58.5719
R1655 VGND.n23 VGND.t13 55.7148
R1656 VGND.n317 VGND.t211 55.7148
R1657 VGND.n310 VGND.t61 55.7148
R1658 VGND.n566 VGND.t22 55.7148
R1659 VGND.n37 VGND.t118 55.7148
R1660 VGND.n38 VGND.t28 55.7148
R1661 VGND.n86 VGND.t40 55.7148
R1662 VGND.n72 VGND.t112 52.8576
R1663 VGND.n153 VGND.t55 52.8576
R1664 VGND.n199 VGND.t5 51.4291
R1665 VGND.n240 VGND.t44 51.4291
R1666 VGND.n23 VGND.t120 40.0005
R1667 VGND.n22 VGND.t9 40.0005
R1668 VGND.n22 VGND.t11 40.0005
R1669 VGND.n346 VGND.t215 40.0005
R1670 VGND.n346 VGND.t209 40.0005
R1671 VGND.n317 VGND.t79 40.0005
R1672 VGND.n112 VGND.t18 40.0005
R1673 VGND.n112 VGND.t20 40.0005
R1674 VGND.n566 VGND.t77 40.0005
R1675 VGND.n37 VGND.t16 40.0005
R1676 VGND.n38 VGND.t3 40.0005
R1677 VGND.n41 VGND.t116 40.0005
R1678 VGND.n41 VGND.t117 40.0005
R1679 VGND.n42 VGND.t32 40.0005
R1680 VGND.n42 VGND.t26 40.0005
R1681 VGND.n82 VGND.t36 40.0005
R1682 VGND.n82 VGND.t38 40.0005
R1683 VGND.n86 VGND.t203 40.0005
R1684 VGND.n645 VGND.t207 38.5719
R1685 VGND.n646 VGND.t58 38.5719
R1686 VGND.n175 VGND.t75 38.5719
R1687 VGND.n174 VGND.t95 38.5719
R1688 VGND.n548 VGND.n547 34.6358
R1689 VGND.n354 VGND.n353 34.6358
R1690 VGND.n355 VGND.n354 34.6358
R1691 VGND.n371 VGND.n369 34.6358
R1692 VGND.n661 VGND.n71 34.6358
R1693 VGND.n71 VGND.n70 34.6358
R1694 VGND.n544 VGND.n543 34.6358
R1695 VGND.n191 VGND.n145 28.8787
R1696 VGND.n199 VGND.t87 28.7917
R1697 VGND.n240 VGND.t83 28.7917
R1698 VGND.n72 VGND.t42 27.5691
R1699 VGND.n153 VGND.t73 27.5691
R1700 VGND.n310 VGND.t71 26.8576
R1701 VGND.n385 VGND.n375 26.6009
R1702 VGND.n168 VGND.n167 25.7355
R1703 VGND.n592 VGND.n575 25.6926
R1704 VGND.n193 VGND.n191 25.6926
R1705 VGND.n347 VGND.n345 25.6005
R1706 VGND.n603 VGND.n113 25.6005
R1707 VGND.n65 VGND.n64 25.6005
R1708 VGND.n503 VGND.t15 25.4291
R1709 VGND.n527 VGND.t205 25.4291
R1710 VGND.n498 VGND.t67 24.9236
R1711 VGND.n498 VGND.t51 24.9236
R1712 VGND.n497 VGND.t47 24.9236
R1713 VGND.n497 VGND.t105 24.9236
R1714 VGND.n530 VGND.t93 24.9236
R1715 VGND.n530 VGND.t103 24.9236
R1716 VGND.n144 VGND.t114 24.9236
R1717 VGND.n144 VGND.t106 24.9236
R1718 VGND.n152 VGND.t89 24.9236
R1719 VGND.n152 VGND.t101 24.9236
R1720 VGND.n658 VGND.n74 24.7086
R1721 VGND.n348 VGND.n347 24.4711
R1722 VGND.n353 VGND.n318 24.4711
R1723 VGND.n565 VGND.n113 24.4711
R1724 VGND.n575 VGND.n574 24.4711
R1725 VGND.n70 VGND.n39 24.4711
R1726 VGND.n66 VGND.n65 24.4711
R1727 VGND.n348 VGND.n318 24.0946
R1728 VGND.n574 VGND.n565 24.0946
R1729 VGND.n66 VGND.n39 24.0946
R1730 VGND.n537 VGND.n532 24.0946
R1731 VGND.n386 VGND.n308 23.7181
R1732 VGND.n386 VGND.n385 23.7181
R1733 VGND.n537 VGND.n536 23.7181
R1734 VGND.n168 VGND.n154 23.7181
R1735 VGND.n73 VGND.t69 22.3257
R1736 VGND.n345 VGND.n320 19.9534
R1737 VGND.n604 VGND.n603 19.9534
R1738 VGND.n64 VGND.n43 19.9534
R1739 VGND.n541 VGND.n532 19.9534
R1740 VGND.n605 VGND.n604 19.914
R1741 VGND.n341 VGND.n320 19.3355
R1742 VGND.n531 VGND.n528 18.4476
R1743 VGND.n526 VGND.n525 18.0316
R1744 VGND.n647 VGND.n644 17.961
R1745 VGND.n176 VGND.n173 17.9321
R1746 VGND.n300 VGND.n299 17.6577
R1747 VGND.n682 VGND.n681 17.3181
R1748 VGND.n60 VGND.n43 17.3181
R1749 VGND.n418 VGND.n417 17.195
R1750 VGND.n172 VGND.n154 16.9417
R1751 VGND.t182 VGND.t37 16.8587
R1752 VGND.n355 VGND.n311 16.1887
R1753 VGND.n450 VGND.n127 16.0722
R1754 VGND.n659 VGND.n658 15.8123
R1755 VGND.n636 VGND.n635 15.6833
R1756 VGND.n660 VGND.n659 15.4358
R1757 VGND.n246 VGND.n245 15.3963
R1758 VGND.n371 VGND.n370 15.0593
R1759 VGND.n585 VGND.n578 14.8179
R1760 VGND.n161 VGND.n160 14.8179
R1761 VGND.n644 VGND.n77 14.775
R1762 VGND.n544 VGND.n531 14.3064
R1763 VGND.n474 VGND.n473 14.2735
R1764 VGND.n681 VGND.n680 11.9186
R1765 VGND.n337 VGND.n336 9.71789
R1766 VGND.n581 VGND.n580 9.71789
R1767 VGND.n474 VGND.n469 9.3005
R1768 VGND.n477 VGND.n476 9.3005
R1769 VGND.n478 VGND.n468 9.3005
R1770 VGND.n480 VGND.n479 9.3005
R1771 VGND.n482 VGND.n123 9.3005
R1772 VGND.n484 VGND.n483 9.3005
R1773 VGND.n467 VGND.n122 9.3005
R1774 VGND.n466 VGND.n465 9.3005
R1775 VGND.n455 VGND.n124 9.3005
R1776 VGND.n454 VGND.n453 9.3005
R1777 VGND.n452 VGND.n126 9.3005
R1778 VGND.n450 VGND.n449 9.3005
R1779 VGND.n682 VGND.n18 9.3005
R1780 VGND.n681 VGND.n10 9.3005
R1781 VGND.n680 VGND.n679 9.3005
R1782 VGND.n678 VGND.n677 9.3005
R1783 VGND.n675 VGND.n21 9.3005
R1784 VGND.n674 VGND.n673 9.3005
R1785 VGND.n672 VGND.n24 9.3005
R1786 VGND.n395 VGND.n25 9.3005
R1787 VGND.n397 VGND.n396 9.3005
R1788 VGND.n407 VGND.n406 9.3005
R1789 VGND.n411 VGND.n410 9.3005
R1790 VGND.n413 VGND.n412 9.3005
R1791 VGND.n415 VGND.n414 9.3005
R1792 VGND.n417 VGND.n416 9.3005
R1793 VGND.n418 VGND.n138 9.3005
R1794 VGND.n421 VGND.n420 9.3005
R1795 VGND.n422 VGND.n137 9.3005
R1796 VGND.n424 VGND.n423 9.3005
R1797 VGND.n426 VGND.n425 9.3005
R1798 VGND.n427 VGND.n131 9.3005
R1799 VGND.n439 VGND.n438 9.3005
R1800 VGND.n441 VGND.n440 9.3005
R1801 VGND.n443 VGND.n442 9.3005
R1802 VGND.n444 VGND.n128 9.3005
R1803 VGND.n447 VGND.n446 9.3005
R1804 VGND.n448 VGND.n127 9.3005
R1805 VGND.n583 VGND.n579 9.3005
R1806 VGND.n586 VGND.n585 9.3005
R1807 VGND.n589 VGND.n588 9.3005
R1808 VGND.n590 VGND.n564 9.3005
R1809 VGND.n593 VGND.n592 9.3005
R1810 VGND.n575 VGND.n563 9.3005
R1811 VGND.n574 VGND.n573 9.3005
R1812 VGND.n565 VGND.n114 9.3005
R1813 VGND.n601 VGND.n113 9.3005
R1814 VGND.n603 VGND.n602 9.3005
R1815 VGND.n604 VGND.n111 9.3005
R1816 VGND.n606 VGND.n605 9.3005
R1817 VGND.n608 VGND.n607 9.3005
R1818 VGND.n609 VGND.n108 9.3005
R1819 VGND.n611 VGND.n610 9.3005
R1820 VGND.n612 VGND.n106 9.3005
R1821 VGND.n620 VGND.n619 9.3005
R1822 VGND.n622 VGND.n621 9.3005
R1823 VGND.n105 VGND.n103 9.3005
R1824 VGND.n379 VGND.n378 9.3005
R1825 VGND.n380 VGND.n376 9.3005
R1826 VGND.n382 VGND.n381 9.3005
R1827 VGND.n383 VGND.n375 9.3005
R1828 VGND.n339 VGND.n321 9.3005
R1829 VGND.n342 VGND.n341 9.3005
R1830 VGND.n343 VGND.n320 9.3005
R1831 VGND.n345 VGND.n344 9.3005
R1832 VGND.n347 VGND.n319 9.3005
R1833 VGND.n349 VGND.n348 9.3005
R1834 VGND.n350 VGND.n318 9.3005
R1835 VGND.n353 VGND.n352 9.3005
R1836 VGND.n354 VGND.n316 9.3005
R1837 VGND.n356 VGND.n355 9.3005
R1838 VGND.n369 VGND.n368 9.3005
R1839 VGND.n372 VGND.n371 9.3005
R1840 VGND.n373 VGND.n308 9.3005
R1841 VGND.n386 VGND.n374 9.3005
R1842 VGND.n385 VGND.n384 9.3005
R1843 VGND.n538 VGND.n537 9.3005
R1844 VGND.n539 VGND.n532 9.3005
R1845 VGND.n541 VGND.n540 9.3005
R1846 VGND.n543 VGND.n529 9.3005
R1847 VGND.n545 VGND.n544 9.3005
R1848 VGND.n547 VGND.n546 9.3005
R1849 VGND.n549 VGND.n548 9.3005
R1850 VGND.n525 VGND.n494 9.3005
R1851 VGND.n523 VGND.n493 9.3005
R1852 VGND.n521 VGND.n520 9.3005
R1853 VGND.n519 VGND.n499 9.3005
R1854 VGND.n518 VGND.n517 9.3005
R1855 VGND.n515 VGND.n500 9.3005
R1856 VGND.n514 VGND.n513 9.3005
R1857 VGND.n512 VGND.n511 9.3005
R1858 VGND.n510 VGND.n502 9.3005
R1859 VGND.n509 VGND.n508 9.3005
R1860 VGND.n506 VGND.n505 9.3005
R1861 VGND.n635 VGND.n634 9.3005
R1862 VGND.n60 VGND.n59 9.3005
R1863 VGND.n62 VGND.n43 9.3005
R1864 VGND.n64 VGND.n63 9.3005
R1865 VGND.n65 VGND.n40 9.3005
R1866 VGND.n67 VGND.n66 9.3005
R1867 VGND.n68 VGND.n39 9.3005
R1868 VGND.n70 VGND.n69 9.3005
R1869 VGND.n71 VGND.n35 9.3005
R1870 VGND.n662 VGND.n661 9.3005
R1871 VGND.n658 VGND.n657 9.3005
R1872 VGND.n650 VGND.n649 9.3005
R1873 VGND.n648 VGND.n76 9.3005
R1874 VGND.n642 VGND.n77 9.3005
R1875 VGND.n641 VGND.n640 9.3005
R1876 VGND.n639 VGND.n79 9.3005
R1877 VGND.n636 VGND.n84 9.3005
R1878 VGND.n644 VGND.n643 9.3005
R1879 VGND.n255 VGND.n233 9.3005
R1880 VGND.n258 VGND.n257 9.3005
R1881 VGND.n237 VGND.n232 9.3005
R1882 VGND.n236 VGND.n235 9.3005
R1883 VGND.n269 VGND.n268 9.3005
R1884 VGND.n270 VGND.n223 9.3005
R1885 VGND.n272 VGND.n271 9.3005
R1886 VGND.n273 VGND.n222 9.3005
R1887 VGND.n252 VGND.n251 9.3005
R1888 VGND.n250 VGND.n238 9.3005
R1889 VGND.n249 VGND.n248 9.3005
R1890 VGND.n246 VGND.n239 9.3005
R1891 VGND.n275 VGND.n274 9.3005
R1892 VGND.n277 VGND.n221 9.3005
R1893 VGND.n279 VGND.n278 9.3005
R1894 VGND.n281 VGND.n280 9.3005
R1895 VGND.n160 VGND.n0 9.3005
R1896 VGND.n161 VGND.n156 9.3005
R1897 VGND.n165 VGND.n164 9.3005
R1898 VGND.n167 VGND.n166 9.3005
R1899 VGND.n169 VGND.n168 9.3005
R1900 VGND.n170 VGND.n154 9.3005
R1901 VGND.n172 VGND.n171 9.3005
R1902 VGND.n177 VGND.n151 9.3005
R1903 VGND.n179 VGND.n178 9.3005
R1904 VGND.n191 VGND.n190 9.3005
R1905 VGND.n194 VGND.n193 9.3005
R1906 VGND.n195 VGND.n141 9.3005
R1907 VGND.n303 VGND.n302 9.3005
R1908 VGND.n301 VGND.n300 9.3005
R1909 VGND.n299 VGND.n298 9.3005
R1910 VGND.n297 VGND.n296 9.3005
R1911 VGND.n295 VGND.n198 9.3005
R1912 VGND.n293 VGND.n292 9.3005
R1913 VGND.n202 VGND.n201 9.3005
R1914 VGND.n216 VGND.n215 9.3005
R1915 VGND.n217 VGND.n206 9.3005
R1916 VGND.n284 VGND.n283 9.3005
R1917 VGND.n649 VGND.n648 9.05896
R1918 VGND.n178 VGND.n177 9.05896
R1919 VGND.n548 VGND.n526 8.28285
R1920 VGND.n675 VGND.n674 8.23546
R1921 VGND.n674 VGND.n24 8.23546
R1922 VGND.n395 VGND.n24 8.23546
R1923 VGND.n381 VGND.n380 8.23546
R1924 VGND.n380 VGND.n379 8.23546
R1925 VGND.n379 VGND.n105 8.23546
R1926 VGND.n621 VGND.n105 8.23546
R1927 VGND.n621 VGND.n620 8.23546
R1928 VGND.n620 VGND.n106 8.23546
R1929 VGND.n610 VGND.n609 8.23546
R1930 VGND.n609 VGND.n608 8.23546
R1931 VGND.n510 VGND.n509 8.23546
R1932 VGND.n511 VGND.n510 8.23546
R1933 VGND.n515 VGND.n514 8.23546
R1934 VGND.n517 VGND.n515 8.23546
R1935 VGND.n521 VGND.n499 8.23546
R1936 VGND.n296 VGND.n295 8.23546
R1937 VGND.n252 VGND.n238 8.23546
R1938 VGND.n676 VGND.n675 8.05644
R1939 VGND.n294 VGND.n293 8.05644
R1940 VGND.n543 VGND.n542 7.90638
R1941 VGND.n509 VGND.n504 7.78791
R1942 VGND.n511 VGND.n501 7.78791
R1943 VGND.n677 VGND.n20 7.6984
R1944 VGND.n414 VGND.n139 7.6984
R1945 VGND.n381 VGND.n377 7.6984
R1946 VGND.n608 VGND.n110 7.6984
R1947 VGND.n505 VGND.n87 7.6984
R1948 VGND.n522 VGND.n521 7.6984
R1949 VGND.n524 VGND.n523 7.6984
R1950 VGND.n248 VGND.n247 7.6984
R1951 VGND.n296 VGND.n200 7.60889
R1952 VGND.n241 VGND.n238 7.60889
R1953 VGND.n396 VGND.n395 6.88949
R1954 VGND.n414 VGND.n413 6.88949
R1955 VGND.n293 VGND.n201 6.88949
R1956 VGND.n173 VGND.n172 6.77697
R1957 VGND.n590 VGND.n589 6.26433
R1958 VGND.n640 VGND.n639 6.26433
R1959 VGND.n303 VGND.n141 6.26433
R1960 VGND.n275 VGND.n222 6.02861
R1961 VGND.n340 VGND.n339 5.98311
R1962 VGND.n584 VGND.n583 5.98311
R1963 VGND.n164 VGND.n162 5.98311
R1964 VGND.n591 VGND.n590 5.85582
R1965 VGND.n192 VGND.n141 5.85582
R1966 VGND.n640 VGND.n81 5.51539
R1967 VGND.n542 VGND.n541 5.27109
R1968 VGND.n682 VGND.n11 5.13108
R1969 VGND.n682 VGND.n19 5.13108
R1970 VGND.n473 VGND.n470 5.13108
R1971 VGND.n473 VGND.n471 5.13108
R1972 VGND.n60 VGND.n45 5.13108
R1973 VGND.n60 VGND.n46 5.13108
R1974 VGND.n536 VGND.n533 5.13108
R1975 VGND.n536 VGND.n534 5.13108
R1976 VGND.n160 VGND.n157 5.13108
R1977 VGND.n160 VGND.n159 5.13108
R1978 VGND.n245 VGND.n242 5.13108
R1979 VGND.n245 VGND.n244 5.13108
R1980 VGND.n339 VGND.n338 4.8005
R1981 VGND.n583 VGND.n582 4.8005
R1982 VGND.n164 VGND.n163 4.8005
R1983 VGND.n420 VGND.n137 4.67352
R1984 VGND.n424 VGND.n137 4.67352
R1985 VGND.n425 VGND.n424 4.67352
R1986 VGND.n425 VGND.n131 4.67352
R1987 VGND.n439 VGND.n131 4.67352
R1988 VGND.n440 VGND.n439 4.67352
R1989 VGND.n444 VGND.n443 4.67352
R1990 VGND.n446 VGND.n444 4.67352
R1991 VGND.n453 VGND.n452 4.67352
R1992 VGND.n453 VGND.n124 4.67352
R1993 VGND.n466 VGND.n124 4.67352
R1994 VGND.n467 VGND.n466 4.67352
R1995 VGND.n483 VGND.n467 4.67352
R1996 VGND.n483 VGND.n482 4.67352
R1997 VGND.n480 VGND.n468 4.67352
R1998 VGND.n476 VGND.n468 4.67352
R1999 VGND.n278 VGND.n277 4.67352
R2000 VGND.n271 VGND.n270 4.67352
R2001 VGND.n270 VGND.n269 4.67352
R2002 VGND.n237 VGND.n236 4.67352
R2003 VGND.n257 VGND.n237 4.67352
R2004 VGND.n683 VGND.n682 4.62124
R2005 VGND.n61 VGND.n60 4.62124
R2006 VGND.n636 VGND.n85 4.62124
R2007 VGND.n160 VGND.n158 4.62124
R2008 VGND.n182 VGND.n150 4.51401
R2009 VGND.n187 VGND.n143 4.51401
R2010 VGND.n430 VGND.n136 4.51401
R2011 VGND.n435 VGND.n130 4.51401
R2012 VGND.n696 VGND.n1 4.51401
R2013 VGND.n56 VGND.n44 4.51401
R2014 VGND.n333 VGND.n323 4.51401
R2015 VGND.n685 VGND.n684 4.51401
R2016 VGND.n228 VGND.n226 4.51401
R2017 VGND.n260 VGND.n259 4.51401
R2018 VGND.n558 VGND.n491 4.51401
R2019 VGND.n496 VGND.n495 4.51401
R2020 VGND.n600 VGND.n599 4.51401
R2021 VGND.n595 VGND.n594 4.51401
R2022 VGND.n457 VGND.n456 4.51401
R2023 VGND.n486 VGND.n485 4.51401
R2024 VGND.n671 VGND.n670 4.51401
R2025 VGND.n403 VGND.n392 4.51401
R2026 VGND.n665 VGND.n33 4.51401
R2027 VGND.n656 VGND.n655 4.51401
R2028 VGND.n351 VGND.n315 4.51401
R2029 VGND.n365 VGND.n309 4.51401
R2030 VGND.n625 VGND.n101 4.51401
R2031 VGND.n618 VGND.n617 4.51401
R2032 VGND.n97 VGND.n95 4.51401
R2033 VGND.n507 VGND.n93 4.51401
R2034 VGND.n291 VGND.n290 4.51401
R2035 VGND.n286 VGND.n285 4.51401
R2036 VGND.n458 VGND.n125 4.5005
R2037 VGND.n463 VGND.n462 4.5005
R2038 VGND.n464 VGND.n121 4.5005
R2039 VGND.n17 VGND.n16 4.5005
R2040 VGND.n9 VGND.n8 4.5005
R2041 VGND.n429 VGND.n428 4.5005
R2042 VGND.n134 VGND.n132 4.5005
R2043 VGND.n437 VGND.n436 4.5005
R2044 VGND.n394 VGND.n26 4.5005
R2045 VGND.n400 VGND.n398 4.5005
R2046 VGND.n405 VGND.n404 4.5005
R2047 VGND.n567 VGND.n115 4.5005
R2048 VGND.n571 VGND.n570 4.5005
R2049 VGND.n572 VGND.n562 4.5005
R2050 VGND.n327 VGND.n322 4.5005
R2051 VGND.n335 VGND.n334 4.5005
R2052 VGND.n358 VGND.n357 4.5005
R2053 VGND.n359 VGND.n312 4.5005
R2054 VGND.n367 VGND.n366 4.5005
R2055 VGND.n624 VGND.n623 4.5005
R2056 VGND.n613 VGND.n104 4.5005
R2057 VGND.n616 VGND.n107 4.5005
R2058 VGND.n633 VGND.n632 4.5005
R2059 VGND.n91 VGND.n89 4.5005
R2060 VGND.n557 VGND.n556 4.5005
R2061 VGND.n555 VGND.n554 4.5005
R2062 VGND.n551 VGND.n550 4.5005
R2063 VGND.n49 VGND.n47 4.5005
R2064 VGND.n58 VGND.n57 4.5005
R2065 VGND.n664 VGND.n663 4.5005
R2066 VGND.n651 VGND.n36 4.5005
R2067 VGND.n654 VGND.n75 4.5005
R2068 VGND.n96 VGND.n88 4.5005
R2069 VGND.n267 VGND.n266 4.5005
R2070 VGND.n229 VGND.n227 4.5005
R2071 VGND.n234 VGND.n231 4.5005
R2072 VGND.n690 VGND.n689 4.5005
R2073 VGND.n698 VGND.n697 4.5005
R2074 VGND.n181 VGND.n180 4.5005
R2075 VGND.n148 VGND.n146 4.5005
R2076 VGND.n189 VGND.n188 4.5005
R2077 VGND.n210 VGND.n208 4.5005
R2078 VGND.n214 VGND.n213 4.5005
R2079 VGND.n209 VGND.n205 4.5005
R2080 VGND.n420 VGND.n419 4.36875
R2081 VGND.n446 VGND.n445 4.36875
R2082 VGND.n452 VGND.n451 4.36875
R2083 VGND.n476 VGND.n475 4.36875
R2084 VGND.n278 VGND.n220 4.36875
R2085 VGND.n277 VGND.n276 4.36875
R2086 VGND.n271 VGND.n224 4.36875
R2087 VGND.n257 VGND.n256 4.36875
R2088 VGND.n589 VGND.n577 4.28986
R2089 VGND.n638 VGND.n637 4.15369
R2090 VGND.n109 VGND.n106 4.11798
R2091 VGND.n610 VGND.n109 4.11798
R2092 VGND.n517 VGND.n516 4.11798
R2093 VGND.n516 VGND.n499 4.11798
R2094 VGND.n578 VGND.n577 4.07323
R2095 VGND.n637 VGND.n636 4.07323
R2096 VGND.n217 VGND.n216 3.96548
R2097 VGND.n254 VGND.n253 3.79556
R2098 VGND.n407 VGND.n393 3.7069
R2099 VGND.n216 VGND.n207 3.7069
R2100 VGND.n330 VGND.n329 3.48706
R2101 VGND.n52 VGND.n51 3.48706
R2102 VGND.n693 VGND.n692 3.48706
R2103 VGND.n12 VGND.n5 3.45831
R2104 VGND.n287 VGND.n286 3.43925
R2105 VGND.n187 VGND.n186 3.43925
R2106 VGND.n183 VGND.n182 3.43925
R2107 VGND.n435 VGND.n434 3.43925
R2108 VGND.n431 VGND.n430 3.43925
R2109 VGND.n696 VGND.n695 3.43925
R2110 VGND.n56 VGND.n55 3.43925
R2111 VGND.n333 VGND.n332 3.43925
R2112 VGND.n261 VGND.n260 3.43925
R2113 VGND.n263 VGND.n228 3.43925
R2114 VGND.n495 VGND.n489 3.43925
R2115 VGND.n559 VGND.n558 3.43925
R2116 VGND.n596 VGND.n595 3.43925
R2117 VGND.n599 VGND.n598 3.43925
R2118 VGND.n403 VGND.n29 3.43925
R2119 VGND.n670 VGND.n669 3.43925
R2120 VGND.n655 VGND.n30 3.43925
R2121 VGND.n666 VGND.n665 3.43925
R2122 VGND.n617 VGND.n99 3.43925
R2123 VGND.n626 VGND.n625 3.43925
R2124 VGND.n290 VGND.n289 3.43925
R2125 VGND.n629 VGND.n93 3.43925
R2126 VGND.n98 VGND.n97 3.43925
R2127 VGND.n184 VGND.n149 3.4105
R2128 VGND.n185 VGND.n147 3.4105
R2129 VGND.n432 VGND.n135 3.4105
R2130 VGND.n433 VGND.n133 3.4105
R2131 VGND.n691 VGND.n688 3.4105
R2132 VGND.n3 VGND.n2 3.4105
R2133 VGND.n53 VGND.n50 3.4105
R2134 VGND.n54 VGND.n48 3.4105
R2135 VGND.n328 VGND.n326 3.4105
R2136 VGND.n325 VGND.n324 3.4105
R2137 VGND.n687 VGND.n686 3.4105
R2138 VGND.n687 VGND.n5 3.4105
R2139 VGND.n686 VGND.n685 3.4105
R2140 VGND.n14 VGND.n13 3.4105
R2141 VGND.n15 VGND.n7 3.4105
R2142 VGND.n265 VGND.n264 3.4105
R2143 VGND.n262 VGND.n230 3.4105
R2144 VGND.n492 VGND.n490 3.4105
R2145 VGND.n553 VGND.n552 3.4105
R2146 VGND.n568 VGND.n116 3.4105
R2147 VGND.n569 VGND.n561 3.4105
R2148 VGND.n488 VGND.n487 3.4105
R2149 VGND.n488 VGND.n119 3.4105
R2150 VGND.n487 VGND.n486 3.4105
R2151 VGND.n457 VGND.n119 3.4105
R2152 VGND.n460 VGND.n459 3.4105
R2153 VGND.n461 VGND.n120 3.4105
R2154 VGND.n399 VGND.n27 3.4105
R2155 VGND.n402 VGND.n401 3.4105
R2156 VGND.n34 VGND.n32 3.4105
R2157 VGND.n653 VGND.n652 3.4105
R2158 VGND.n364 VGND.n31 3.4105
R2159 VGND.n314 VGND.n31 3.4105
R2160 VGND.n365 VGND.n364 3.4105
R2161 VGND.n315 VGND.n314 3.4105
R2162 VGND.n361 VGND.n360 3.4105
R2163 VGND.n363 VGND.n313 3.4105
R2164 VGND.n102 VGND.n100 3.4105
R2165 VGND.n615 VGND.n614 3.4105
R2166 VGND.n631 VGND.n630 3.4105
R2167 VGND.n92 VGND.n90 3.4105
R2168 VGND.n211 VGND.n203 3.4105
R2169 VGND.n212 VGND.n204 3.4105
R2170 VGND.n661 VGND.n660 3.38874
R2171 VGND.n303 VGND.n142 3.13241
R2172 VGND.n255 VGND.n254 3.05276
R2173 VGND.n473 VGND.n472 3.04861
R2174 VGND.n587 VGND.n578 3.04861
R2175 VGND.n536 VGND.n535 3.04861
R2176 VGND.n245 VGND.n243 3.04861
R2177 VGND.n196 VGND.n142 2.7239
R2178 VGND.n440 VGND.n129 2.33701
R2179 VGND.n443 VGND.n129 2.33701
R2180 VGND.n482 VGND.n481 2.33701
R2181 VGND.n481 VGND.n480 2.33701
R2182 VGND.n269 VGND.n225 2.33701
R2183 VGND.n236 VGND.n225 2.33701
R2184 VGND.n17 VGND.n12 2.33488
R2185 VGND.n329 VGND.n322 2.33488
R2186 VGND.n51 VGND.n47 2.33488
R2187 VGND.n692 VGND.n689 2.33488
R2188 VGND.n369 VGND.n311 2.25932
R2189 VGND.n408 VGND.n407 1.98299
R2190 VGND.n410 VGND.n408 1.98299
R2191 VGND.n410 VGND.n409 1.98299
R2192 VGND.n218 VGND.n217 1.98299
R2193 VGND.n547 VGND.n528 1.88285
R2194 VGND.n409 VGND.n391 1.72441
R2195 VGND.n219 VGND.n218 1.72441
R2196 VGND.n332 VGND.n331 1.69188
R2197 VGND.n331 VGND.n330 1.69188
R2198 VGND.n55 VGND.n6 1.69188
R2199 VGND.n52 VGND.n6 1.69188
R2200 VGND.n695 VGND.n694 1.69188
R2201 VGND.n694 VGND.n693 1.69188
R2202 VGND.n687 VGND.n4 1.69188
R2203 VGND.n597 VGND.n596 1.69188
R2204 VGND.n598 VGND.n597 1.69188
R2205 VGND.n560 VGND.n489 1.69188
R2206 VGND.n560 VGND.n559 1.69188
R2207 VGND.n261 VGND.n117 1.69188
R2208 VGND.n263 VGND.n117 1.69188
R2209 VGND.n488 VGND.n118 1.69188
R2210 VGND.n667 VGND.n30 1.69188
R2211 VGND.n667 VGND.n666 1.69188
R2212 VGND.n668 VGND.n29 1.69188
R2213 VGND.n669 VGND.n668 1.69188
R2214 VGND.n186 VGND.n28 1.69188
R2215 VGND.n183 VGND.n28 1.69188
R2216 VGND.n362 VGND.n31 1.69188
R2217 VGND.n627 VGND.n99 1.69188
R2218 VGND.n627 VGND.n626 1.69188
R2219 VGND.n434 VGND.n94 1.69188
R2220 VGND.n431 VGND.n94 1.69188
R2221 VGND.n288 VGND.n287 1.69188
R2222 VGND.n289 VGND.n288 1.69188
R2223 VGND.n629 VGND.n628 1.69188
R2224 VGND.n628 VGND.n98 1.69188
R2225 VGND.n370 VGND.n308 1.50638
R2226 VGND.n282 VGND.n281 1.40924
R2227 VGND.n283 VGND.n282 1.26145
R2228 VGND.n338 VGND.n337 1.18311
R2229 VGND.n582 VGND.n581 1.18311
R2230 VGND.n163 VGND.n155 1.18311
R2231 VGND.n577 VGND.n576 0.952566
R2232 VGND.n637 VGND.n83 0.952566
R2233 VGND.n248 VGND.n241 0.627073
R2234 VGND.n680 VGND.n20 0.537563
R2235 VGND.n417 VGND.n139 0.537563
R2236 VGND.n377 VGND.n375 0.537563
R2237 VGND.n605 VGND.n110 0.537563
R2238 VGND.n635 VGND.n87 0.537563
R2239 VGND.n523 VGND.n522 0.537563
R2240 VGND.n525 VGND.n524 0.537563
R2241 VGND.n299 VGND.n197 0.537563
R2242 VGND.n247 VGND.n246 0.537563
R2243 VGND.n505 VGND.n504 0.448052
R2244 VGND.n514 VGND.n501 0.448052
R2245 VGND.n341 VGND.n340 0.417891
R2246 VGND.n585 VGND.n584 0.417891
R2247 VGND.n162 VGND.n161 0.417891
R2248 VGND.n167 VGND.n155 0.417891
R2249 VGND.n592 VGND.n591 0.409011
R2250 VGND.n80 VGND.n77 0.409011
R2251 VGND.n193 VGND.n192 0.409011
R2252 VGND.n300 VGND.n196 0.409011
R2253 VGND.n81 VGND.n80 0.340926
R2254 VGND.n419 VGND.n418 0.305262
R2255 VGND.n445 VGND.n127 0.305262
R2256 VGND.n451 VGND.n450 0.305262
R2257 VGND.n475 VGND.n474 0.305262
R2258 VGND.n281 VGND.n220 0.305262
R2259 VGND.n276 VGND.n275 0.305262
R2260 VGND.n224 VGND.n222 0.305262
R2261 VGND.n256 VGND.n255 0.305262
R2262 VGND.n396 VGND.n393 0.259086
R2263 VGND.n413 VGND.n391 0.259086
R2264 VGND.n207 VGND.n201 0.259086
R2265 VGND.n283 VGND.n219 0.259086
R2266 VGND.n588 VGND.n587 0.239726
R2267 VGND.n472 VGND 0.217246
R2268 VGND.n243 VGND 0.217246
R2269 VGND.n535 VGND 0.205527
R2270 VGND.n649 VGND.n74 0.197423
R2271 VGND.n648 VGND.n647 0.197423
R2272 VGND.n177 VGND.n176 0.197423
R2273 VGND.n178 VGND.n145 0.197423
R2274 VGND.n683 VGND.n10 0.180304
R2275 VGND.n62 VGND.n61 0.180304
R2276 VGND.n85 VGND.n79 0.180304
R2277 VGND.n158 VGND.n156 0.180304
R2278 VGND.n677 VGND.n676 0.179521
R2279 VGND.n295 VGND.n294 0.179521
R2280 VGND.n253 VGND.n252 0.179521
R2281 VGND.n694 VGND.n687 0.1603
R2282 VGND.n687 VGND.n6 0.1603
R2283 VGND.n331 VGND.n6 0.1603
R2284 VGND.n488 VGND.n117 0.1603
R2285 VGND.n560 VGND.n488 0.1603
R2286 VGND.n597 VGND.n560 0.1603
R2287 VGND.n668 VGND.n28 0.1603
R2288 VGND.n668 VGND.n667 0.1603
R2289 VGND.n667 VGND.n31 0.1603
R2290 VGND.n288 VGND.n94 0.1603
R2291 VGND.n628 VGND.n94 0.1603
R2292 VGND.n628 VGND.n627 0.1603
R2293 VGND.n472 VGND 0.14207
R2294 VGND.n535 VGND 0.14207
R2295 VGND.n243 VGND 0.14207
R2296 VGND.n587 VGND 0.141725
R2297 VGND.n639 VGND.n638 0.13667
R2298 VGND.n95 VGND.n85 0.134731
R2299 VGND.n679 VGND.n678 0.120292
R2300 VGND.n678 VGND.n21 0.120292
R2301 VGND.n673 VGND.n21 0.120292
R2302 VGND.n673 VGND.n672 0.120292
R2303 VGND.n412 VGND.n411 0.120292
R2304 VGND.n421 VGND.n138 0.120292
R2305 VGND.n422 VGND.n421 0.120292
R2306 VGND.n423 VGND.n422 0.120292
R2307 VGND.n442 VGND.n441 0.120292
R2308 VGND.n442 VGND.n128 0.120292
R2309 VGND.n447 VGND.n128 0.120292
R2310 VGND.n448 VGND.n447 0.120292
R2311 VGND.n449 VGND.n126 0.120292
R2312 VGND.n454 VGND.n126 0.120292
R2313 VGND.n484 VGND.n123 0.120292
R2314 VGND.n479 VGND.n123 0.120292
R2315 VGND.n479 VGND.n478 0.120292
R2316 VGND.n478 VGND.n477 0.120292
R2317 VGND.n477 VGND.n469 0.120292
R2318 VGND.n342 VGND.n321 0.120292
R2319 VGND.n343 VGND.n342 0.120292
R2320 VGND.n344 VGND.n343 0.120292
R2321 VGND.n344 VGND.n319 0.120292
R2322 VGND.n349 VGND.n319 0.120292
R2323 VGND.n350 VGND.n349 0.120292
R2324 VGND.n352 VGND.n350 0.120292
R2325 VGND.n373 VGND.n372 0.120292
R2326 VGND.n383 VGND.n382 0.120292
R2327 VGND.n382 VGND.n376 0.120292
R2328 VGND.n378 VGND.n376 0.120292
R2329 VGND.n612 VGND.n611 0.120292
R2330 VGND.n611 VGND.n108 0.120292
R2331 VGND.n607 VGND.n108 0.120292
R2332 VGND.n607 VGND.n606 0.120292
R2333 VGND.n602 VGND.n111 0.120292
R2334 VGND.n602 VGND.n601 0.120292
R2335 VGND.n593 VGND.n564 0.120292
R2336 VGND.n588 VGND.n564 0.120292
R2337 VGND.n586 VGND.n579 0.120292
R2338 VGND.n580 VGND.n579 0.120292
R2339 VGND.n63 VGND.n62 0.120292
R2340 VGND.n63 VGND.n40 0.120292
R2341 VGND.n67 VGND.n40 0.120292
R2342 VGND.n68 VGND.n67 0.120292
R2343 VGND.n69 VGND.n68 0.120292
R2344 VGND.n650 VGND.n76 0.120292
R2345 VGND.n642 VGND.n641 0.120292
R2346 VGND.n641 VGND.n79 0.120292
R2347 VGND.n508 VGND.n502 0.120292
R2348 VGND.n512 VGND.n502 0.120292
R2349 VGND.n513 VGND.n512 0.120292
R2350 VGND.n518 VGND.n500 0.120292
R2351 VGND.n546 VGND.n545 0.120292
R2352 VGND.n545 VGND.n529 0.120292
R2353 VGND.n540 VGND.n529 0.120292
R2354 VGND.n540 VGND.n539 0.120292
R2355 VGND.n165 VGND.n156 0.120292
R2356 VGND.n166 VGND.n165 0.120292
R2357 VGND.n170 VGND.n169 0.120292
R2358 VGND.n171 VGND.n170 0.120292
R2359 VGND.n195 VGND.n194 0.120292
R2360 VGND.n298 VGND.n297 0.120292
R2361 VGND.n297 VGND.n198 0.120292
R2362 VGND.n292 VGND.n198 0.120292
R2363 VGND.n280 VGND.n279 0.120292
R2364 VGND.n279 VGND.n221 0.120292
R2365 VGND.n274 VGND.n221 0.120292
R2366 VGND.n273 VGND.n272 0.120292
R2367 VGND.n272 VGND.n223 0.120292
R2368 VGND.n258 VGND.n233 0.120292
R2369 VGND.n251 VGND.n250 0.120292
R2370 VGND.n250 VGND.n249 0.120292
R2371 VGND.n249 VGND.n239 0.120292
R2372 VGND.n171 VGND.n150 0.104667
R2373 VGND.n485 VGND.n484 0.102062
R2374 VGND.n546 VGND.n496 0.102062
R2375 VGND.n259 VGND.n258 0.102062
R2376 VGND.n415 VGND 0.0981562
R2377 VGND.n449 VGND 0.0981562
R2378 VGND.n374 VGND 0.0981562
R2379 VGND.n111 VGND 0.0981562
R2380 VGND VGND.n593 0.0981562
R2381 VGND VGND.n586 0.0981562
R2382 VGND.n643 VGND 0.0981562
R2383 VGND VGND.n500 0.0981562
R2384 VGND VGND.n538 0.0981562
R2385 VGND.n169 VGND 0.0981562
R2386 VGND.n298 VGND 0.0981562
R2387 VGND.n280 VGND 0.0981562
R2388 VGND VGND.n273 0.0981562
R2389 VGND.n251 VGND 0.0981562
R2390 VGND.n520 VGND 0.0968542
R2391 VGND.n182 VGND.n181 0.0950946
R2392 VGND.n188 VGND.n187 0.0950946
R2393 VGND.n430 VGND.n429 0.0950946
R2394 VGND.n436 VGND.n435 0.0950946
R2395 VGND.n697 VGND.n696 0.0950946
R2396 VGND.n57 VGND.n56 0.0950946
R2397 VGND.n334 VGND.n333 0.0950946
R2398 VGND.n685 VGND.n8 0.0950946
R2399 VGND.n266 VGND.n228 0.0950946
R2400 VGND.n260 VGND.n231 0.0950946
R2401 VGND.n558 VGND.n557 0.0950946
R2402 VGND.n551 VGND.n495 0.0950946
R2403 VGND.n599 VGND.n115 0.0950946
R2404 VGND.n595 VGND.n562 0.0950946
R2405 VGND.n458 VGND.n457 0.0950946
R2406 VGND.n486 VGND.n121 0.0950946
R2407 VGND.n670 VGND.n26 0.0950946
R2408 VGND.n404 VGND.n403 0.0950946
R2409 VGND.n665 VGND.n664 0.0950946
R2410 VGND.n655 VGND.n654 0.0950946
R2411 VGND.n358 VGND.n315 0.0950946
R2412 VGND.n366 VGND.n365 0.0950946
R2413 VGND.n625 VGND.n624 0.0950946
R2414 VGND.n617 VGND.n616 0.0950946
R2415 VGND.n97 VGND.n96 0.0950946
R2416 VGND.n93 VGND.n91 0.0950946
R2417 VGND.n286 VGND.n205 0.0950946
R2418 VGND.n200 VGND.n197 0.0900105
R2419 VGND.n679 VGND 0.0890417
R2420 VGND VGND.n138 0.0890417
R2421 VGND VGND.n383 0.0890417
R2422 VGND.n692 VGND.n691 0.0878527
R2423 VGND.n51 VGND.n50 0.0878527
R2424 VGND.n329 VGND.n328 0.0878527
R2425 VGND.n14 VGND.n12 0.0878527
R2426 VGND.n416 VGND 0.0877396
R2427 VGND.n384 VGND 0.0877396
R2428 VGND VGND.n642 0.0877396
R2429 VGND VGND.n301 0.0877396
R2430 VGND.n519 VGND 0.0864375
R2431 VGND.n302 VGND 0.0864375
R2432 VGND.n684 VGND.n9 0.0838333
R2433 VGND.n405 VGND.n398 0.0838333
R2434 VGND.n437 VGND.n132 0.0838333
R2435 VGND.n463 VGND.n125 0.0838333
R2436 VGND.n335 VGND.n323 0.0838333
R2437 VGND.n367 VGND.n312 0.0838333
R2438 VGND.n107 VGND.n104 0.0838333
R2439 VGND.n571 VGND.n567 0.0838333
R2440 VGND.n58 VGND.n44 0.0838333
R2441 VGND.n75 VGND.n36 0.0838333
R2442 VGND.n633 VGND.n89 0.0838333
R2443 VGND.n556 VGND.n555 0.0838333
R2444 VGND.n698 VGND.n1 0.0838333
R2445 VGND.n189 VGND.n146 0.0838333
R2446 VGND.n214 VGND.n209 0.0838333
R2447 VGND.n267 VGND.n227 0.0838333
R2448 VGND VGND.n671 0.0825312
R2449 VGND.n428 VGND.n427 0.0825312
R2450 VGND VGND.n351 0.0825312
R2451 VGND.n623 VGND.n622 0.0825312
R2452 VGND VGND.n33 0.0825312
R2453 VGND.n634 VGND.n88 0.0825312
R2454 VGND.n215 VGND.n208 0.0825312
R2455 VGND.n406 VGND.n392 0.078625
R2456 VGND.n368 VGND.n309 0.078625
R2457 VGND.n657 VGND.n656 0.078625
R2458 VGND.n456 VGND.n455 0.0760208
R2459 VGND.n600 VGND.n114 0.0760208
R2460 VGND.n493 VGND.n491 0.0760208
R2461 VGND.n268 VGND.n226 0.0760208
R2462 VGND.n423 VGND.n136 0.0747188
R2463 VGND.n378 VGND.n101 0.0747188
R2464 VGND.n684 VGND.n683 0.0722313
R2465 VGND.n61 VGND.n44 0.0722313
R2466 VGND.n158 VGND.n1 0.0722313
R2467 VGND.n441 VGND.n130 0.0721146
R2468 VGND.n618 VGND.n612 0.0721146
R2469 VGND.n508 VGND.n507 0.0721146
R2470 VGND.n285 VGND.n284 0.0721146
R2471 VGND.n357 VGND.n316 0.0682083
R2472 VGND.n663 VGND.n35 0.0682083
R2473 VGND.n180 VGND.n151 0.0682083
R2474 VGND.n149 VGND.n148 0.0680676
R2475 VGND.n148 VGND.n147 0.0680676
R2476 VGND.n135 VGND.n134 0.0680676
R2477 VGND.n134 VGND.n133 0.0680676
R2478 VGND.n691 VGND.n690 0.0680676
R2479 VGND.n690 VGND.n2 0.0680676
R2480 VGND.n50 VGND.n49 0.0680676
R2481 VGND.n49 VGND.n48 0.0680676
R2482 VGND.n328 VGND.n327 0.0680676
R2483 VGND.n327 VGND.n324 0.0680676
R2484 VGND.n16 VGND.n14 0.0680676
R2485 VGND.n16 VGND.n15 0.0680676
R2486 VGND.n265 VGND.n229 0.0680676
R2487 VGND.n230 VGND.n229 0.0680676
R2488 VGND.n554 VGND.n492 0.0680676
R2489 VGND.n554 VGND.n553 0.0680676
R2490 VGND.n570 VGND.n568 0.0680676
R2491 VGND.n570 VGND.n569 0.0680676
R2492 VGND.n462 VGND.n460 0.0680676
R2493 VGND.n462 VGND.n461 0.0680676
R2494 VGND.n400 VGND.n399 0.0680676
R2495 VGND.n402 VGND.n400 0.0680676
R2496 VGND.n651 VGND.n34 0.0680676
R2497 VGND.n653 VGND.n651 0.0680676
R2498 VGND.n360 VGND.n359 0.0680676
R2499 VGND.n359 VGND.n313 0.0680676
R2500 VGND.n613 VGND.n102 0.0680676
R2501 VGND.n615 VGND.n613 0.0680676
R2502 VGND.n632 VGND.n90 0.0680676
R2503 VGND.n632 VGND.n631 0.0680676
R2504 VGND.n290 VGND 0.0680676
R2505 VGND.n213 VGND.n211 0.0680676
R2506 VGND.n213 VGND.n212 0.0680676
R2507 VGND.n464 VGND.n122 0.0656042
R2508 VGND.n572 VGND.n563 0.0656042
R2509 VGND.n550 VGND.n549 0.0656042
R2510 VGND.n234 VGND.n232 0.0656042
R2511 VGND.n18 VGND.n17 0.0590938
R2512 VGND.n336 VGND.n322 0.0590938
R2513 VGND.n59 VGND.n47 0.0590938
R2514 VGND.n689 VGND.n0 0.0590938
R2515 VGND VGND.n143 0.0577917
R2516 VGND.n204 VGND.n203 0.0574697
R2517 VGND.n185 VGND.n184 0.0574697
R2518 VGND.n433 VGND.n432 0.0574697
R2519 VGND.n688 VGND.n3 0.0574697
R2520 VGND.n54 VGND.n53 0.0574697
R2521 VGND.n326 VGND.n325 0.0574697
R2522 VGND.n13 VGND.n5 0.0574697
R2523 VGND.n686 VGND.n7 0.0574697
R2524 VGND.n264 VGND.n262 0.0574697
R2525 VGND.n552 VGND.n490 0.0574697
R2526 VGND.n561 VGND.n116 0.0574697
R2527 VGND.n459 VGND.n119 0.0574697
R2528 VGND.n487 VGND.n120 0.0574697
R2529 VGND.n401 VGND.n27 0.0574697
R2530 VGND.n652 VGND.n32 0.0574697
R2531 VGND.n361 VGND.n314 0.0574697
R2532 VGND.n364 VGND.n363 0.0574697
R2533 VGND.n614 VGND.n100 0.0574697
R2534 VGND.n630 VGND.n92 0.0574697
R2535 VGND.n465 VGND.n464 0.0551875
R2536 VGND.n573 VGND.n572 0.0551875
R2537 VGND.n235 VGND.n234 0.0551875
R2538 VGND.n397 VGND.n394 0.0525833
R2539 VGND.n357 VGND.n356 0.0525833
R2540 VGND.n663 VGND.n662 0.0525833
R2541 VGND.n180 VGND.n179 0.0525833
R2542 VGND.n438 VGND.n130 0.0486771
R2543 VGND.n619 VGND.n618 0.0486771
R2544 VGND.n507 VGND.n506 0.0486771
R2545 VGND.n285 VGND.n206 0.0486771
R2546 VGND.n426 VGND.n136 0.0460729
R2547 VGND.n103 VGND.n101 0.0460729
R2548 VGND.n95 VGND.n84 0.0460729
R2549 VGND.n291 VGND.n202 0.0460729
R2550 VGND.n456 VGND.n454 0.0447708
R2551 VGND.n601 VGND.n600 0.0447708
R2552 VGND.n520 VGND.n491 0.0447708
R2553 VGND.n226 VGND.n223 0.0447708
R2554 VGND VGND.n291 0.0434688
R2555 VGND.n411 VGND.n392 0.0421667
R2556 VGND.n372 VGND.n309 0.0421667
R2557 VGND.n656 VGND.n650 0.0421667
R2558 VGND.n194 VGND.n143 0.0421667
R2559 VGND.n181 VGND.n149 0.0410405
R2560 VGND.n188 VGND.n147 0.0410405
R2561 VGND.n429 VGND.n135 0.0410405
R2562 VGND.n436 VGND.n133 0.0410405
R2563 VGND.n697 VGND.n2 0.0410405
R2564 VGND.n57 VGND.n48 0.0410405
R2565 VGND.n334 VGND.n324 0.0410405
R2566 VGND.n15 VGND.n8 0.0410405
R2567 VGND.n266 VGND.n265 0.0410405
R2568 VGND.n231 VGND.n230 0.0410405
R2569 VGND.n557 VGND.n492 0.0410405
R2570 VGND.n553 VGND.n551 0.0410405
R2571 VGND.n568 VGND.n115 0.0410405
R2572 VGND.n569 VGND.n562 0.0410405
R2573 VGND.n460 VGND.n458 0.0410405
R2574 VGND.n461 VGND.n121 0.0410405
R2575 VGND.n399 VGND.n26 0.0410405
R2576 VGND.n404 VGND.n402 0.0410405
R2577 VGND.n664 VGND.n34 0.0410405
R2578 VGND.n654 VGND.n653 0.0410405
R2579 VGND.n360 VGND.n358 0.0410405
R2580 VGND.n366 VGND.n313 0.0410405
R2581 VGND.n624 VGND.n102 0.0410405
R2582 VGND.n616 VGND.n615 0.0410405
R2583 VGND.n96 VGND.n90 0.0410405
R2584 VGND.n631 VGND.n91 0.0410405
R2585 VGND.n211 VGND.n210 0.0410405
R2586 VGND.n212 VGND.n205 0.0410405
R2587 VGND.n428 VGND.n426 0.0382604
R2588 VGND.n623 VGND.n103 0.0382604
R2589 VGND.n208 VGND.n202 0.0382604
R2590 VGND.n394 VGND 0.0369583
R2591 VGND.n438 VGND.n437 0.0356562
R2592 VGND.n619 VGND.n107 0.0356562
R2593 VGND.n506 VGND.n89 0.0356562
R2594 VGND.n209 VGND.n206 0.0356562
R2595 VGND VGND.n518 0.0343542
R2596 VGND VGND.n195 0.0343542
R2597 VGND VGND.n415 0.0330521
R2598 VGND VGND.n374 0.0330521
R2599 VGND.n550 VGND 0.0330521
R2600 VGND.n302 VGND 0.0330521
R2601 VGND VGND.n10 0.03175
R2602 VGND VGND.n25 0.03175
R2603 VGND.n398 VGND.n397 0.03175
R2604 VGND.n356 VGND.n312 0.03175
R2605 VGND.n384 VGND 0.03175
R2606 VGND.n662 VGND.n36 0.03175
R2607 VGND.n538 VGND 0.03175
R2608 VGND.n179 VGND.n146 0.03175
R2609 VGND.n292 VGND 0.03175
R2610 VGND.n289 VGND.n203 0.0292489
R2611 VGND.n330 VGND.n326 0.0292489
R2612 VGND.n332 VGND.n325 0.0292489
R2613 VGND.n53 VGND.n52 0.0292489
R2614 VGND.n55 VGND.n54 0.0292489
R2615 VGND.n693 VGND.n688 0.0292489
R2616 VGND.n695 VGND.n3 0.0292489
R2617 VGND.n7 VGND.n4 0.0292489
R2618 VGND.n13 VGND.n4 0.0292489
R2619 VGND.n598 VGND.n116 0.0292489
R2620 VGND.n596 VGND.n561 0.0292489
R2621 VGND.n559 VGND.n490 0.0292489
R2622 VGND.n552 VGND.n489 0.0292489
R2623 VGND.n264 VGND.n263 0.0292489
R2624 VGND.n262 VGND.n261 0.0292489
R2625 VGND.n120 VGND.n118 0.0292489
R2626 VGND.n459 VGND.n118 0.0292489
R2627 VGND.n666 VGND.n32 0.0292489
R2628 VGND.n652 VGND.n30 0.0292489
R2629 VGND.n669 VGND.n27 0.0292489
R2630 VGND.n401 VGND.n29 0.0292489
R2631 VGND.n184 VGND.n183 0.0292489
R2632 VGND.n186 VGND.n185 0.0292489
R2633 VGND.n363 VGND.n362 0.0292489
R2634 VGND.n362 VGND.n361 0.0292489
R2635 VGND.n626 VGND.n100 0.0292489
R2636 VGND.n614 VGND.n99 0.0292489
R2637 VGND.n432 VGND.n431 0.0292489
R2638 VGND.n434 VGND.n433 0.0292489
R2639 VGND.n287 VGND.n204 0.0292489
R2640 VGND.n98 VGND.n92 0.0292489
R2641 VGND.n630 VGND.n629 0.0292489
R2642 VGND.n465 VGND.n463 0.0291458
R2643 VGND.n573 VGND.n571 0.0291458
R2644 VGND.n555 VGND.n494 0.0291458
R2645 VGND.n235 VGND.n227 0.0291458
R2646 VGND.n210 VGND 0.027527
R2647 VGND VGND.n519 0.0239375
R2648 VGND.n18 VGND 0.0226354
R2649 VGND.n672 VGND 0.0226354
R2650 VGND.n412 VGND 0.0226354
R2651 VGND.n416 VGND 0.0226354
R2652 VGND VGND.n448 0.0226354
R2653 VGND VGND.n469 0.0226354
R2654 VGND.n336 VGND 0.0226354
R2655 VGND.n352 VGND 0.0226354
R2656 VGND VGND.n373 0.0226354
R2657 VGND.n606 VGND 0.0226354
R2658 VGND.n580 VGND 0.0226354
R2659 VGND.n59 VGND 0.0226354
R2660 VGND.n69 VGND 0.0226354
R2661 VGND VGND.n76 0.0226354
R2662 VGND VGND.n84 0.0226354
R2663 VGND.n513 VGND 0.0226354
R2664 VGND VGND.n494 0.0226354
R2665 VGND.n539 VGND 0.0226354
R2666 VGND VGND.n0 0.0226354
R2667 VGND.n166 VGND 0.0226354
R2668 VGND.n301 VGND 0.0226354
R2669 VGND.n284 VGND 0.0226354
R2670 VGND.n274 VGND 0.0226354
R2671 VGND VGND.n233 0.0226354
R2672 VGND VGND.n239 0.0226354
R2673 VGND.n643 VGND 0.0213333
R2674 VGND.n190 VGND 0.0213333
R2675 VGND.n485 VGND.n122 0.0187292
R2676 VGND.n594 VGND.n563 0.0187292
R2677 VGND.n549 VGND.n496 0.0187292
R2678 VGND.n259 VGND.n232 0.0187292
R2679 VGND.n671 VGND.n25 0.016125
R2680 VGND.n351 VGND.n316 0.016125
R2681 VGND.n35 VGND.n33 0.016125
R2682 VGND.n88 VGND 0.016125
R2683 VGND.n151 VGND.n150 0.016125
R2684 VGND.n323 VGND.n321 0.0122188
R2685 VGND.n455 VGND.n125 0.0083125
R2686 VGND.n567 VGND.n114 0.0083125
R2687 VGND.n556 VGND.n493 0.0083125
R2688 VGND.n268 VGND.n267 0.0083125
R2689 VGND.n331 VGND 0.00755
R2690 VGND.n597 VGND 0.00755
R2691 VGND.n31 VGND 0.00755
R2692 VGND.n627 VGND 0.00755
R2693 VGND.n406 VGND.n405 0.00570833
R2694 VGND.n368 VGND.n367 0.00570833
R2695 VGND.n657 VGND.n75 0.00570833
R2696 VGND.n190 VGND.n189 0.00570833
R2697 VGND.n594 VGND 0.00440625
R2698 VGND VGND.n9 0.00310417
R2699 VGND VGND.n335 0.00310417
R2700 VGND VGND.n58 0.00310417
R2701 VGND VGND.n698 0.00310417
R2702 VGND.n427 VGND.n132 0.00180208
R2703 VGND.n622 VGND.n104 0.00180208
R2704 VGND.n634 VGND.n633 0.00180208
R2705 VGND.n215 VGND.n214 0.00180208
R2706 n[0].n9 n[0].n8 332.332
R2707 n[0].n9 n[0].n7 296.493
R2708 n[0].n2 n[0].n0 135.248
R2709 n[0].n6 n[0].n5 98.982
R2710 n[0].n2 n[0].n1 98.981
R2711 n[0].n4 n[0].n3 98.981
R2712 n[0].n11 n[0].n6 42.0805
R2713 n[0].n4 n[0].n2 36.2672
R2714 n[0].n6 n[0].n4 36.2672
R2715 n[0].n7 n[0].t8 26.5955
R2716 n[0].n7 n[0].t10 26.5955
R2717 n[0].n8 n[0].t9 26.5955
R2718 n[0].n8 n[0].t11 26.5955
R2719 n[0] n[0].n11 26.0019
R2720 n[0].n0 n[0].t2 24.9236
R2721 n[0].n0 n[0].t3 24.9236
R2722 n[0].n1 n[0].t1 24.9236
R2723 n[0].n1 n[0].t0 24.9236
R2724 n[0].n3 n[0].t7 24.9236
R2725 n[0].n3 n[0].t5 24.9236
R2726 n[0].n5 n[0].t6 24.9236
R2727 n[0].n5 n[0].t4 24.9236
R2728 n[0].n10 n[0].n9 18.5605
R2729 n[0].n11 n[0].n10 2.0805
R2730 n[0].n10 n[0] 0.6405
R2731 n[1].n3 n[1].n1 647.148
R2732 n[1].n6 n[1].n0 243.627
R2733 n[1].n3 n[1].n2 194.441
R2734 n[1].n8 n[1].n7 185
R2735 n[1].n7 n[1].t3 40.0005
R2736 n[1].n7 n[1].t0 40.0005
R2737 n[1].n0 n[1].t1 40.0005
R2738 n[1].n0 n[1].t2 40.0005
R2739 n[1].n2 n[1].t7 27.5805
R2740 n[1].n2 n[1].t4 27.5805
R2741 n[1].n1 n[1].t5 27.5805
R2742 n[1].n1 n[1].t6 27.5805
R2743 n[1] n[1].n8 24.248
R2744 n[1] n[1].n4 19.2609
R2745 n[1].n4 n[1].n3 15.5262
R2746 n[1].n8 n[1].n6 15.262
R2747 n[1].n5 n[1] 9.00791
R2748 n[1].n6 n[1].n5 6.77697
R2749 n[1].n4 n[1] 2.70819
R2750 n[1].n5 n[1] 1.73877
R2751 p[3].n6 p[3].n5 256.104
R2752 p[3].n9 p[3].n7 243.68
R2753 p[3].n2 p[3].n0 241.847
R2754 p[3].n9 p[3].n8 205.28
R2755 p[3].n6 p[3].n4 202.094
R2756 p[3].n2 p[3].n1 185
R2757 p[3].n4 p[3].t5 26.5955
R2758 p[3].n4 p[3].t7 26.5955
R2759 p[3].n7 p[3].t10 26.5955
R2760 p[3].n7 p[3].t9 26.5955
R2761 p[3].n8 p[3].t11 26.5955
R2762 p[3].n8 p[3].t8 26.5955
R2763 p[3].n5 p[3].t6 26.5955
R2764 p[3].n5 p[3].t4 26.5955
R2765 p[3].n1 p[3].t2 24.9236
R2766 p[3].n1 p[3].t0 24.9236
R2767 p[3].n0 p[3].t3 24.9236
R2768 p[3].n0 p[3].t1 24.9236
R2769 p[3] p[3].n9 22.9652
R2770 p[3].n3 p[3].n2 20.9279
R2771 p[3].n3 p[3] 15.3283
R2772 p[3].n10 p[3].n6 13.9299
R2773 p[3].n10 p[3] 13.9299
R2774 p[3] p[3].n10 5.26405
R2775 p[3].n10 p[3] 2.87153
R2776 p[3] p[3].n3 2.03414
R2777 n[3].n2 n[3].n0 647.148
R2778 n[3].n6 n[3].n4 243.627
R2779 n[3].n6 n[3].n5 200.262
R2780 n[3].n2 n[3].n1 194.441
R2781 n[3].n4 n[3].t0 40.0005
R2782 n[3].n4 n[3].t1 40.0005
R2783 n[3].n5 n[3].t2 40.0005
R2784 n[3].n5 n[3].t3 40.0005
R2785 n[3].n1 n[3].t6 27.5805
R2786 n[3].n1 n[3].t7 27.5805
R2787 n[3].n0 n[3].t4 27.5805
R2788 n[3].n0 n[3].t5 27.5805
R2789 n[3] n[3].n8 23.4037
R2790 n[3] n[3].n3 19.2609
R2791 n[3].n3 n[3].n2 15.5262
R2792 n[3].n8 n[3] 8.05976
R2793 n[3].n7 n[3].n6 6.77697
R2794 n[3].n3 n[3] 2.70819
R2795 n[3].n7 n[3] 1.73877
R2796 n[3].n8 n[3].n7 0.948648
R2797 p[1].n5 p[1].n4 647.148
R2798 p[1].n2 p[1].n0 243.627
R2799 p[1].n2 p[1].n1 200.262
R2800 p[1].n5 p[1].n3 194.441
R2801 p[1].n0 p[1].t0 40.0005
R2802 p[1].n0 p[1].t1 40.0005
R2803 p[1].n1 p[1].t2 40.0005
R2804 p[1].n1 p[1].t3 40.0005
R2805 p[1].n3 p[1].t4 27.5805
R2806 p[1].n3 p[1].t5 27.5805
R2807 p[1].n4 p[1].t6 27.5805
R2808 p[1].n4 p[1].t7 27.5805
R2809 p[1] p[1].n6 17.2864
R2810 p[1] p[1].n2 10.4115
R2811 p[1] p[1].n5 9.86463
R2812 p[1].n6 p[1] 8.05976
R2813 p[1].n6 p[1] 2.68692
R2814 n[2].n5 n[2].n4 647.148
R2815 n[2].n2 n[2].n0 243.627
R2816 n[2].n2 n[2].n1 200.262
R2817 n[2].n5 n[2].n3 194.441
R2818 n[2].n0 n[2].t2 40.0005
R2819 n[2].n0 n[2].t3 40.0005
R2820 n[2].n1 n[2].t0 40.0005
R2821 n[2].n1 n[2].t1 40.0005
R2822 n[2].n3 n[2].t5 27.5805
R2823 n[2].n3 n[2].t6 27.5805
R2824 n[2].n4 n[2].t7 27.5805
R2825 n[2].n4 n[2].t4 27.5805
R2826 n[2] n[2].n6 24.7742
R2827 n[2].n6 n[2] 15.365
R2828 n[2] n[2].n2 10.4115
R2829 n[2] n[2].n5 9.86463
R2830 n[2].n6 n[2] 4.18512
R2831 p[2].n1 p[2].n0 642.239
R2832 p[2].n8 p[2].n7 585
R2833 p[2].n9 p[2].n8 290.56
R2834 p[2].n4 p[2].n2 243.627
R2835 p[2].n4 p[2].n3 200.262
R2836 p[2].n2 p[2].t2 40.0005
R2837 p[2].n2 p[2].t3 40.0005
R2838 p[2].n3 p[2].t0 40.0005
R2839 p[2].n3 p[2].t1 40.0005
R2840 p[2].n8 p[2].t4 27.5805
R2841 p[2].n8 p[2].t5 27.5805
R2842 p[2].n0 p[2].t6 27.5805
R2843 p[2].n0 p[2].t7 27.5805
R2844 p[2].n6 p[2] 19.2609
R2845 p[2] p[2].n9 15.9794
R2846 p[2].n7 p[2].n1 14.7697
R2847 p[2] p[2].n5 9.00791
R2848 p[2].n9 p[2].n1 8.03728
R2849 p[2].n5 p[2].n4 6.77697
R2850 p[2].n7 p[2].n6 5.90819
R2851 p[2].n6 p[2] 2.70819
R2852 p[2].n5 p[2] 1.73877
R2853 p[0].n2 p[0].n0 647.148
R2854 p[0].n6 p[0].n4 243.627
R2855 p[0].n6 p[0].n5 200.262
R2856 p[0].n2 p[0].n1 194.441
R2857 p[0].n4 p[0].t2 40.0005
R2858 p[0].n4 p[0].t3 40.0005
R2859 p[0].n5 p[0].t0 40.0005
R2860 p[0].n5 p[0].t1 40.0005
R2861 p[0] p[0].n8 33.1212
R2862 p[0].n1 p[0].t4 27.5805
R2863 p[0].n1 p[0].t5 27.5805
R2864 p[0].n0 p[0].t6 27.5805
R2865 p[0].n0 p[0].t7 27.5805
R2866 p[0] p[0].n3 19.2609
R2867 p[0].n3 p[0].n2 15.5262
R2868 p[0].n8 p[0] 8.05976
R2869 p[0].n7 p[0].n6 6.77697
R2870 p[0].n3 p[0] 2.70819
R2871 p[0].n7 p[0] 1.73877
R2872 p[0].n8 p[0].n7 0.948648
R2873 a.n0 a.t1 276.464
R2874 a.n0 a.t0 196.131
R2875 a.n1 a.n0 153.385
R2876 a.n1 a 10.0713
R2877 a a.n1 2.94104
R2878 b.n0 b.t1 276.464
R2879 b.n0 b.t0 196.131
R2880 b.n1 b.n0 152
R2881 b.n1 b 10.783
R2882 b b.n1 1.55726
C0 p[0] a_5179_2767# 0.001818f
C1 a_2599_3677# VPWR 0.190042f
C2 _01_ net1 0.183603f
C3 a_4842_2473# net1 9.5e-19
C4 net1 n[0] 0.680517f
C5 net2 a_3523_2767# 0.239365f
C6 a_4903_5263# a_5179_4399# 1.67e-19
C7 net2 p[3] 0.557656f
C8 n[1] a_2879_2223# 0.336811f
C9 a_5179_2767# _04_ 0.422447f
C10 net1 n[3] 1.17e-19
C11 a_4760_2473# a_4819_2883# 0.001329f
C12 n[1] _00_ 0.020945f
C13 net2 a_5177_5737# 0.002523f
C14 a_5179_2767# a_5179_3311# 0.052341f
C15 net1 a_5179_2767# 0.001824f
C16 a_5095_5737# p[3] 0.017866f
C17 net1 a_2879_2223# 0.002006f
C18 p[1] a_4075_2767# 5.17e-19
C19 net1 _00_ 0.096879f
C20 a_4627_3127# VPWR 0.080484f
C21 VPWR p[2] 0.874521f
C22 a_5179_2223# p[1] 8.94e-19
C23 a_3703_2767# a_4075_2767# 0.001895f
C24 a_5177_5737# a_5095_5737# 0.005162f
C25 VPWR a_5179_4399# 0.556376f
C26 net2 b 0.380065f
C27 n[2] _02_ 9.03e-19
C28 net2 p[1] 0.00218f
C29 net2 a_4075_2767# 0.082281f
C30 a_4760_2473# _03_ 0.10634f
C31 net1 a_2419_3677# 0.223081f
C32 net1 a_2327_5487# 0.201662f
C33 a_5179_2223# net2 9.56e-19
C34 a_3703_2767# net2 0.064477f
C35 b a_5095_5737# 0.052438f
C36 n[1] n[2] 0.02803f
C37 n[2] _04_ 0.006062f
C38 a_2557_2767# n[1] 9.65e-19
C39 a_4627_3127# a_4819_2883# 0.101254f
C40 net1 n[2] 0.568369f
C41 a_3793_3133# VPWR 4.34e-19
C42 a_2557_2767# net1 0.181933f
C43 a_4903_5493# a_4903_5263# 4.2e-19
C44 net2 a_5095_5737# 0.152191f
C45 _01_ n[0] 6.9e-20
C46 net1 a_4903_5263# 0.218905f
C47 _02_ VPWR 0.355242f
C48 p[0] VPWR 0.549795f
C49 a_4627_3127# a_4901_2883# 3.5e-20
C50 _01_ a_5179_2767# 1.09e-20
C51 a_4751_3339# VPWR 0.217067f
C52 a_5179_2223# a_4760_2473# 0.001f
C53 _03_ a_5179_4399# 4.58e-20
C54 _01_ _00_ 9.69e-19
C55 n[0] _00_ 0.041057f
C56 p[3] p[2] 0.002059f
C57 VPWR a_4903_5493# 0.078375f
C58 n[1] VPWR 0.367301f
C59 VPWR _04_ 0.157277f
C60 net2 a_4760_2473# 0.171637f
C61 p[3] a_5179_4399# 0.003762f
C62 VPWR a_5179_3311# 0.437791f
C63 n[3] a_5179_2767# 8.94e-19
C64 net1 VPWR 4.08889f
C65 n[0] a_2419_3677# 0.00168f
C66 net1 a 0.060808f
C67 a_2879_2223# _00_ 0.25164f
C68 _05_ a_4903_5263# 0.01603f
C69 _02_ a_4819_2883# 0.009399f
C70 a_2599_3677# a_2689_3311# 0.004764f
C71 net2 a_2599_3677# 0.203551f
C72 a_4627_3127# p[1] 6.03e-19
C73 a_4751_3339# a_4819_2883# 0.003659f
C74 b p[2] 3.51e-20
C75 a_4627_3127# a_4075_2767# 0.001493f
C76 p[1] p[2] 3.35e-19
C77 _01_ n[2] 0.02282f
C78 a_4312_5461# a_4903_5493# 0.002785f
C79 a_2419_3677# _00_ 0.001633f
C80 a_4819_2883# _04_ 0.121744f
C81 a_2557_2767# _01_ 3.44e-19
C82 a_2557_2767# n[0] 0.255994f
C83 _03_ _02_ 0.410893f
C84 _02_ a_4901_2883# 7.28e-20
C85 net1 a_4819_2883# 0.136683f
C86 net1 a_4312_5461# 0.05084f
C87 _05_ VPWR 0.513343f
C88 p[0] _03_ 0.031468f
C89 a_4627_3127# net2 0.186914f
C90 n[3] n[2] 0.001766f
C91 net2 p[2] 0.006494f
C92 a_4751_3339# _03_ 0.01704f
C93 n[2] a_5179_2767# 6.56e-20
C94 a_2879_2223# n[2] 6.55e-19
C95 net2 a_5179_4399# 0.014558f
C96 n[2] _00_ 3.49e-19
C97 a_2557_2767# a_2879_2223# 0.001238f
C98 _03_ a_4837_3339# 7.44e-20
C99 a_2557_2767# _00_ 0.026107f
C100 _03_ _04_ 0.1429f
C101 a_4901_2883# _04_ 3.82e-19
C102 _03_ a_5179_3311# 0.203359f
C103 net1 _03_ 0.020464f
C104 a_4903_5493# p[3] 0.008402f
C105 net1 a_4901_2883# 0.001856f
C106 net1 a_3523_2767# 0.137644f
C107 a_5179_3311# p[3] 2.13e-20
C108 net1 p[3] 0.225569f
C109 _01_ VPWR 0.141427f
C110 a_4842_2473# VPWR 0.002134f
C111 n[0] VPWR 0.352414f
C112 a_3703_2767# a_3793_3133# 0.004764f
C113 a_2557_2767# a_2419_3677# 1.07e-19
C114 a_5177_5737# a_4903_5493# 3.5e-20
C115 a_4312_5461# _05_ 2.96e-19
C116 p[1] _02_ 9.94e-19
C117 a_4075_2767# _02_ 1.21e-21
C118 net2 a_3793_3133# 0.001719f
C119 p[0] p[1] 0.067253f
C120 n[3] VPWR 0.52858f
C121 a_5179_2223# _02_ 0.246074f
C122 VPWR a_5179_2767# 0.422804f
C123 a_2879_2223# VPWR 0.496359f
C124 a_5179_2223# p[0] 8.93e-19
C125 b a_4903_5493# 0.039708f
C126 VPWR _00_ 0.492287f
C127 a_2557_2767# n[2] 1.15e-19
C128 net2 _02_ 0.119334f
C129 p[1] _04_ 0.023051f
C130 a_4075_2767# _04_ 2.18e-19
C131 net1 b 0.191923f
C132 _03_ _05_ 1.32e-19
C133 net2 p[0] 0.002127f
C134 p[1] a_5179_3311# 9.86e-19
C135 net1 p[1] 0.001109f
C136 net1 a_4075_2767# 0.072889f
C137 _01_ a_4819_2883# 3.36e-20
C138 a_5179_2223# _04_ 1.11e-19
C139 net2 a_4751_3339# 0.097252f
C140 _05_ p[3] 0.239496f
C141 a_2419_3677# VPWR 0.260273f
C142 a_3703_2767# net1 0.233026f
C143 net2 a_4903_5493# 0.123859f
C144 net2 n[1] 5.85e-19
C145 net2 a_4837_3339# 9.11e-19
C146 a_2327_5487# VPWR 0.369627f
C147 net2 _04_ 0.012497f
C148 net1 a_2689_3311# 5.55e-19
C149 net2 a_5179_3311# 0.00588f
C150 net2 net1 1.45741f
C151 a_5177_5737# _05_ 7.86e-19
C152 a_5179_2767# a_4819_2883# 0.002083f
C153 a_2327_5487# a 0.173221f
C154 a_5095_5737# a_4903_5493# 0.101254f
C155 a_4842_2473# _03_ 4.96e-19
C156 n[2] VPWR 0.570613f
C157 net1 a_5095_5737# 0.00232f
C158 a_2557_2767# VPWR 0.664434f
C159 _01_ a_3523_2767# 0.001089f
C160 a_4760_2473# _02_ 0.018215f
C161 b _05_ 0.075495f
C162 p[2] a_5179_4399# 0.337919f
C163 VPWR a_4903_5263# 0.028248f
C164 n[3] _03_ 0.001259f
C165 _03_ a_5179_2767# 0.050375f
C166 a_4760_2473# a_4751_3339# 4.34e-19
C167 n[1] a_4760_2473# 2.34e-20
C168 net2 _05_ 0.11267f
C169 a_3523_2767# _00_ 0.00183f
C170 net1 a_4760_2473# 0.125892f
C171 n[2] a_4819_2883# 0.009294f
C172 _01_ p[1] 1.37e-19
C173 _01_ a_4075_2767# 0.408145f
C174 _05_ a_5095_5737# 0.123524f
C175 a_3703_2767# _01_ 0.093531f
C176 a VPWR 0.387516f
C177 a_4627_3127# _02_ 4.73e-19
C178 net1 a_2599_3677# 0.014286f
C179 n[3] p[1] 0.00746f
C180 _01_ net2 0.134826f
C181 a_4842_2473# net2 5.11e-19
C182 p[1] a_5179_2767# 0.339173f
C183 a_4075_2767# a_5179_2767# 3.74e-21
C184 net2 n[0] 0.173347f
C185 p[0] p[2] 0.001063f
C186 _02_ a_5179_4399# 2.19e-19
C187 _03_ n[2] 0.004102f
C188 n[2] a_4901_2883# 1.11e-19
C189 a_4627_3127# a_4751_3339# 5.45e-19
C190 a_5179_2223# n[3] 0.329355f
C191 a_4075_2767# _00_ 0.001298f
C192 p[0] a_5179_4399# 1.15e-19
C193 n[2] a_3523_2767# 2.52e-19
C194 a_5179_2223# a_5179_2767# 0.050529f
C195 a_2557_2767# a_3523_2767# 0.01539f
C196 a_4627_3127# _04_ 0.00129f
C197 a_3703_2767# _00_ 0.001845f
C198 net2 n[3] 2.41e-19
C199 net2 a_5179_2767# 0.002254f
C200 a_4627_3127# net1 0.139449f
C201 a_4312_5461# VPWR 0.35757f
C202 VPWR a_4819_2883# 0.123093f
C203 a_2689_3311# _00_ 0.001544f
C204 a_5179_3311# p[2] 5.47e-20
C205 net2 a_2879_2223# 0.036218f
C206 net1 p[2] 0.001016f
C207 p[3] a_4903_5263# 0.189438f
C208 net2 _00_ 0.122695f
C209 a_5179_3311# a_5179_4399# 0.001652f
C210 net1 a_5179_4399# 0.001694f
C211 net2 a_2419_3677# 0.095435f
C212 _03_ VPWR 0.534521f
C213 a_4842_2473# a_4760_2473# 0.004767f
C214 VPWR a_4901_2883# 0.0012f
C215 n[2] p[1] 2.33e-19
C216 n[2] a_4075_2767# 0.33834f
C217 a_3523_2767# VPWR 0.234232f
C218 VPWR p[3] 1.03748f
C219 p[0] _02_ 0.002263f
C220 a_3703_2767# n[2] 3.97e-19
C221 a_5179_2223# n[2] 0.002384f
C222 n[3] a_4760_2473# 1.35e-19
C223 net1 a_3793_3133# 2.66e-19
C224 a_4751_3339# _02_ 0.110488f
C225 _05_ p[2] 0.035813f
C226 net2 n[2] 0.276603f
C227 a_5177_5737# VPWR 6.34e-19
C228 a_2557_2767# net2 0.210178f
C229 n[0] a_2599_3677# 0.001372f
C230 a_4837_3339# _02_ 0.001478f
C231 _05_ a_5179_4399# 0.245904f
C232 _02_ _04_ 0.053416f
C233 _02_ a_5179_3311# 0.203053f
C234 net1 _02_ 0.008948f
C235 net2 a_4903_5263# 0.080227f
C236 p[0] a_5179_3311# 0.329185f
C237 a_4751_3339# a_4837_3339# 0.006584f
C238 net1 p[0] 4.07e-19
C239 _03_ a_4819_2883# 0.002857f
C240 a_4901_2883# a_4819_2883# 0.005162f
C241 b VPWR 0.608191f
C242 a_4751_3339# a_5179_3311# 0.001175f
C243 net1 a_4751_3339# 0.193587f
C244 p[1] VPWR 0.57701f
C245 a_4075_2767# VPWR 0.438039f
C246 a_2599_3677# _00_ 0.084911f
C247 a_5095_5737# a_4903_5263# 4.68e-19
C248 a_4627_3127# _01_ 9.39e-20
C249 a_4312_5461# p[3] 1.52e-19
C250 net1 a_4903_5493# 0.153574f
C251 net1 n[1] 1.33e-19
C252 net1 a_4837_3339# 0.001645f
C253 a_5179_3311# _04_ 4.96e-20
C254 net1 _04_ 0.006601f
C255 a_5179_2223# VPWR 0.423176f
C256 a_3703_2767# VPWR 0.168337f
C257 net1 a_5179_3311# 0.003382f
C258 a_2689_3311# VPWR 0.001077f
C259 net2 VPWR 4.40655f
C260 a_4760_2473# n[2] 0.008879f
C261 a_2419_3677# a_2599_3677# 0.185422f
C262 _03_ p[3] 1.91e-21
C263 _02_ _05_ 0.002132f
C264 VPWR a_5095_5737# 0.12582f
C265 a_4312_5461# b 0.17615f
C266 p[1] a_4819_2883# 4.97e-19
C267 a_4075_2767# a_4819_2883# 0.001003f
C268 _01_ a_3793_3133# 8.17e-20
C269 _05_ a_4903_5493# 0.003327f
C270 a_5177_5737# p[3] 0.00107f
C271 _05_ a_5179_3311# 6.3e-19
C272 net1 _05_ 0.060099f
C273 net2 a_4819_2883# 0.040325f
C274 net2 a_4312_5461# 0.190752f
C275 _01_ _02_ 6.09e-21
C276 _03_ p[1] 0.034297f
C277 a_4760_2473# VPWR 0.180101f
C278 a_4627_3127# n[2] 0.042087f
C279 b p[3] 0.136111f
C280 a_3793_3133# _00_ 1.94e-19
C281 a_4312_5461# a_5095_5737# 1.44e-19
C282 a_5179_2223# _03_ 0.170725f
C283 n[3] _02_ 0.022864f
C284 _02_ a_5179_2767# 0.019263f
C285 a_3703_2767# a_3523_2767# 0.185422f
C286 n[3] p[0] 0.550473f
C287 _01_ _04_ 7.72e-19
C288 net2 _03_ 0.096664f
C289 b a_5177_5737# 9.84e-19
C290 net2 a_4901_2883# 0.001173f
C291 n[3] VGND 1.6058f
C292 n[1] VGND 1.43826f
C293 p[1] VGND 1.58512f
C294 n[2] VGND 1.33075f
C295 n[0] VGND 2.32339f
C296 p[0] VGND 2.131f
C297 p[2] VGND 1.56136f
C298 p[3] VGND 1.69075f
C299 b VGND 1.24771f
C300 a VGND 1.22032f
C301 VPWR VGND 83.42087f
C302 a_4842_2473# VGND 0.001581f
C303 a_5179_2223# VGND 0.570586f
C304 a_4760_2473# VGND 0.26415f
C305 a_2879_2223# VGND 0.68829f
C306 a_4901_2883# VGND 3.42e-19
C307 a_5179_2767# VGND 0.544f
C308 _04_ VGND 0.281424f
C309 a_4819_2883# VGND 0.280043f
C310 a_4627_3127# VGND 0.306654f
C311 a_2557_2767# VGND 0.050875f
C312 a_3793_3133# VGND 0.005478f
C313 a_4075_2767# VGND 0.576904f
C314 _01_ VGND 0.289986f
C315 a_3703_2767# VGND 0.248329f
C316 a_3523_2767# VGND 0.243777f
C317 a_4837_3339# VGND 0.007629f
C318 _02_ VGND 0.661432f
C319 a_2689_3311# VGND 0.005471f
C320 _00_ VGND 0.879193f
C321 a_5179_3311# VGND 0.577895f
C322 _03_ VGND 0.624442f
C323 a_4751_3339# VGND 0.312074f
C324 a_2599_3677# VGND 0.255292f
C325 a_2419_3677# VGND 0.259064f
C326 a_5179_4399# VGND 0.574241f
C327 a_4903_5263# VGND 0.610445f
C328 _05_ VGND 0.72125f
C329 a_5177_5737# VGND 2.26e-19
C330 a_4903_5493# VGND 0.329899f
C331 a_5095_5737# VGND 0.254516f
C332 net2 VGND 4.35326f
C333 net1 VGND 5.46581f
C334 a_4312_5461# VGND 0.351481f
C335 a_2327_5487# VGND 0.350093f
C336 VPWR.t72 VGND 0.002945f
C337 VPWR.n0 VGND 0.007958f
C338 VPWR.n1 VGND 0.003451f
C339 VPWR.t232 VGND 0.006139f
C340 VPWR.t27 VGND 0.002945f
C341 VPWR.n2 VGND 0.001723f
C342 VPWR.n3 VGND 0.001201f
C343 VPWR.n4 VGND 0.001157f
C344 VPWR.n5 VGND 0.002063f
C345 VPWR.n6 VGND 0.001995f
C346 VPWR.n7 VGND 0.001995f
C347 VPWR.n8 VGND 0.136057f
C348 VPWR.n9 VGND 0.002063f
C349 VPWR.n10 VGND 0.001728f
C350 VPWR.n11 VGND 9.25e-19
C351 VPWR.n12 VGND 0.001201f
C352 VPWR.n13 VGND 0.001201f
C353 VPWR.n14 VGND 0.001807f
C354 VPWR.n15 VGND 0.001728f
C355 VPWR.t104 VGND 0.001055f
C356 VPWR.t118 VGND 0.001055f
C357 VPWR.n16 VGND 0.002265f
C358 VPWR.t15 VGND 0.001094f
C359 VPWR.t17 VGND 0.001094f
C360 VPWR.n17 VGND 0.002219f
C361 VPWR.t120 VGND 0.003975f
C362 VPWR.t13 VGND 0.004579f
C363 VPWR.t83 VGND 0.002945f
C364 VPWR.t240 VGND 0.006251f
C365 VPWR.n19 VGND 0.016026f
C366 VPWR.t84 VGND 0.002945f
C367 VPWR.n20 VGND 0.008729f
C368 VPWR.t90 VGND 0.002945f
C369 VPWR.t223 VGND 0.006251f
C370 VPWR.n22 VGND 0.016026f
C371 VPWR.t91 VGND 0.002945f
C372 VPWR.n23 VGND 0.008729f
C373 VPWR.n24 VGND 0.007385f
C374 VPWR.n25 VGND 0.003286f
C375 VPWR.n26 VGND 0.004675f
C376 VPWR.n27 VGND 4.92e-19
C377 VPWR.n28 VGND 0.004318f
C378 VPWR.n29 VGND 0.003754f
C379 VPWR.n30 VGND 8.9e-19
C380 VPWR.n31 VGND 6.24e-19
C381 VPWR.n32 VGND 0.002081f
C382 VPWR.n33 VGND 0.002569f
C383 VPWR.t19 VGND 0.001485f
C384 VPWR.t196 VGND 0.001094f
C385 VPWR.n34 VGND 0.002741f
C386 VPWR.t124 VGND 0.001055f
C387 VPWR.t184 VGND 0.001055f
C388 VPWR.n35 VGND 0.002265f
C389 VPWR.n36 VGND 0.002582f
C390 VPWR.t165 VGND 0.001055f
C391 VPWR.t182 VGND 0.001055f
C392 VPWR.n37 VGND 0.002265f
C393 VPWR.n38 VGND 0.00239f
C394 VPWR.t175 VGND 0.004153f
C395 VPWR.n39 VGND 0.003517f
C396 VPWR.n40 VGND 4.53e-19
C397 VPWR.t226 VGND 0.012382f
C398 VPWR.t10 VGND 0.002921f
C399 VPWR.n41 VGND 0.012258f
C400 VPWR.n42 VGND 0.013485f
C401 VPWR.t11 VGND 0.002965f
C402 VPWR.n43 VGND 0.003466f
C403 VPWR.n44 VGND 4.31e-19
C404 VPWR.t82 VGND 0.034947f
C405 VPWR.t12 VGND 0.031408f
C406 VPWR.t119 VGND 0.009511f
C407 VPWR.t14 VGND 0.00929f
C408 VPWR.t103 VGND 0.009511f
C409 VPWR.t16 VGND 0.00929f
C410 VPWR.t117 VGND 0.009511f
C411 VPWR.t18 VGND 0.00929f
C412 VPWR.t123 VGND 0.010617f
C413 VPWR.t195 VGND 0.00929f
C414 VPWR.t183 VGND 0.007299f
C415 VPWR.t164 VGND 0.009953f
C416 VPWR.t181 VGND 0.013382f
C417 VPWR.t174 VGND 0.016368f
C418 VPWR.t204 VGND 0.02046f
C419 VPWR.t9 VGND 0.008295f
C420 VPWR.t43 VGND 0.030524f
C421 VPWR.t85 VGND 0.122095f
C422 VPWR.t68 VGND 0.122095f
C423 VPWR.n45 VGND 0.018757f
C424 VPWR.t213 VGND 0.003214f
C425 VPWR.t69 VGND 0.003214f
C426 VPWR.n46 VGND 0.004383f
C427 VPWR.n47 VGND 0.001276f
C428 VPWR.n48 VGND 0.001201f
C429 VPWR.n49 VGND 9.25e-19
C430 VPWR.n50 VGND 0.001728f
C431 VPWR.n51 VGND 0.002063f
C432 VPWR.n52 VGND 0.074031f
C433 VPWR.n54 VGND 0.002012f
C434 VPWR.n55 VGND 0.105044f
C435 VPWR.n56 VGND 0.002063f
C436 VPWR.n57 VGND 0.001157f
C437 VPWR.n58 VGND 0.001201f
C438 VPWR.n59 VGND 0.003451f
C439 VPWR.t225 VGND 0.016877f
C440 VPWR.n60 VGND 0.007399f
C441 VPWR.n61 VGND 0.007027f
C442 VPWR.n62 VGND 0.00179f
C443 VPWR.t54 VGND 0.030303f
C444 VPWR.t187 VGND 0.014156f
C445 VPWR.t189 VGND 0.019022f
C446 VPWR.t191 VGND 0.019022f
C447 VPWR.t193 VGND 0.020128f
C448 VPWR.t33 VGND 0.017916f
C449 VPWR.t23 VGND 0.018469f
C450 VPWR.t129 VGND 0.017031f
C451 VPWR.t172 VGND 0.021234f
C452 VPWR.t109 VGND 0.02046f
C453 VPWR.t6 VGND 0.030524f
C454 VPWR.t168 VGND 0.018027f
C455 VPWR.t0 VGND 0.02057f
C456 VPWR.t115 VGND 0.029418f
C457 VPWR.t199 VGND 0.019907f
C458 VPWR.t49 VGND 0.013603f
C459 VPWR.t147 VGND 0.05784f
C460 VPWR.t215 VGND 0.064255f
C461 VPWR.t57 VGND 0.050873f
C462 VPWR.n63 VGND 0.02215f
C463 VPWR.n64 VGND 0.003097f
C464 VPWR.n65 VGND 0.003451f
C465 VPWR.t173 VGND 8.87e-19
C466 VPWR.t130 VGND 3.31e-19
C467 VPWR.n66 VGND 0.004047f
C468 VPWR.n67 VGND 0.00435f
C469 VPWR.n68 VGND 0.002983f
C470 VPWR.t218 VGND 0.04257f
C471 VPWR.t194 VGND 0.001485f
C472 VPWR.t34 VGND 0.001094f
C473 VPWR.n69 VGND 0.002741f
C474 VPWR.t190 VGND 0.001094f
C475 VPWR.t192 VGND 0.001094f
C476 VPWR.n70 VGND 0.002219f
C477 VPWR.n71 VGND 0.003978f
C478 VPWR.n72 VGND 0.001726f
C479 VPWR.n73 VGND 0.001157f
C480 VPWR.n74 VGND 0.002063f
C481 VPWR.n75 VGND 9.25e-19
C482 VPWR.n76 VGND 0.001519f
C483 VPWR.t188 VGND 0.004625f
C484 VPWR.n77 VGND 0.005361f
C485 VPWR.t55 VGND 0.002945f
C486 VPWR.t230 VGND 0.006251f
C487 VPWR.n79 VGND 0.016026f
C488 VPWR.t56 VGND 0.002945f
C489 VPWR.n80 VGND 0.008729f
C490 VPWR.t97 VGND 0.002945f
C491 VPWR.t247 VGND 0.006251f
C492 VPWR.n82 VGND 0.016026f
C493 VPWR.t98 VGND 0.002945f
C494 VPWR.n83 VGND 0.008729f
C495 VPWR.n84 VGND 0.007265f
C496 VPWR.n85 VGND 0.003286f
C497 VPWR.n86 VGND 0.004281f
C498 VPWR.n87 VGND 0.001157f
C499 VPWR.n88 VGND 0.001995f
C500 VPWR.n89 VGND 0.001807f
C501 VPWR.n90 VGND 0.001278f
C502 VPWR.n91 VGND 0.001201f
C503 VPWR.n92 VGND 0.001434f
C504 VPWR.t24 VGND 0.003214f
C505 VPWR.n93 VGND 0.002497f
C506 VPWR.n94 VGND 0.002081f
C507 VPWR.n95 VGND 0.001201f
C508 VPWR.n96 VGND 0.001407f
C509 VPWR.n97 VGND 0.001157f
C510 VPWR.n98 VGND 9.25e-19
C511 VPWR.n99 VGND 0.002063f
C512 VPWR.n100 VGND 0.001995f
C513 VPWR.n101 VGND 0.001807f
C514 VPWR.n102 VGND 0.001728f
C515 VPWR.n103 VGND 0.001201f
C516 VPWR.n104 VGND 0.004161f
C517 VPWR.n105 VGND 0.00589f
C518 VPWR.n106 VGND 0.0013f
C519 VPWR.n107 VGND 0.019884f
C520 VPWR.n108 VGND 0.003192f
C521 VPWR.n109 VGND 0.002045f
C522 VPWR.n110 VGND 0.003133f
C523 VPWR.n111 VGND 0.003451f
C524 VPWR.n112 VGND 0.003168f
C525 VPWR.n113 VGND 0.005832f
C526 VPWR.n114 VGND 0.003357f
C527 VPWR.t110 VGND 0.00177f
C528 VPWR.n115 VGND 0.005176f
C529 VPWR.n116 VGND 0.003428f
C530 VPWR.n117 VGND 0.003451f
C531 VPWR.n118 VGND 0.002045f
C532 VPWR.n119 VGND 4.53e-19
C533 VPWR.n120 VGND 0.00182f
C534 VPWR.n121 VGND 0.00947f
C535 VPWR.t25 VGND 0.003226f
C536 VPWR.n122 VGND 0.003669f
C537 VPWR.t58 VGND 0.002942f
C538 VPWR.n123 VGND 0.001367f
C539 VPWR.n124 VGND 0.002128f
C540 VPWR.n125 VGND 4.31e-19
C541 VPWR.n126 VGND 0.001276f
C542 VPWR.n127 VGND 0.001157f
C543 VPWR.n128 VGND 0.002063f
C544 VPWR.n129 VGND 9.25e-19
C545 VPWR.n130 VGND 9.25e-19
C546 VPWR.n131 VGND 0.001157f
C547 VPWR.n132 VGND 0.001407f
C548 VPWR.n133 VGND 0.001726f
C549 VPWR.n134 VGND 0.001201f
C550 VPWR.n135 VGND 0.005979f
C551 VPWR.t216 VGND 0.003214f
C552 VPWR.n136 VGND 0.003435f
C553 VPWR.n137 VGND 0.010605f
C554 VPWR.n138 VGND 0.009075f
C555 VPWR.t229 VGND 0.04257f
C556 VPWR.n139 VGND 0.003289f
C557 VPWR.n140 VGND 0.003451f
C558 VPWR.t148 VGND 0.003214f
C559 VPWR.n141 VGND 0.004061f
C560 VPWR.t237 VGND 0.04257f
C561 VPWR.n142 VGND 0.021448f
C562 VPWR.n143 VGND 0.001201f
C563 VPWR.n144 VGND 0.001157f
C564 VPWR.n145 VGND 0.002063f
C565 VPWR.n146 VGND 0.136057f
C566 VPWR.n147 VGND 0.001995f
C567 VPWR.n148 VGND 0.001995f
C568 VPWR.n149 VGND 0.002063f
C569 VPWR.n150 VGND 0.001728f
C570 VPWR.n151 VGND 9.25e-19
C571 VPWR.n152 VGND 0.001201f
C572 VPWR.t3 VGND 6.73e-19
C573 VPWR.t114 VGND 4.43e-19
C574 VPWR.n153 VGND 0.001149f
C575 VPWR.n154 VGND 0.003647f
C576 VPWR.n155 VGND 0.003133f
C577 VPWR.t235 VGND 0.04257f
C578 VPWR.n156 VGND 0.019884f
C579 VPWR.n157 VGND 0.003414f
C580 VPWR.t75 VGND 0.001485f
C581 VPWR.t198 VGND 0.001094f
C582 VPWR.n158 VGND 0.002741f
C583 VPWR.t79 VGND 0.001094f
C584 VPWR.t81 VGND 0.001094f
C585 VPWR.n159 VGND 0.002219f
C586 VPWR.t145 VGND 0.003214f
C587 VPWR.n160 VGND 0.002497f
C588 VPWR.n161 VGND 0.001726f
C589 VPWR.n162 VGND 0.001157f
C590 VPWR.n163 VGND 0.002063f
C591 VPWR.n164 VGND 9.25e-19
C592 VPWR.t106 VGND 0.0018f
C593 VPWR.t141 VGND 0.034947f
C594 VPWR.t60 VGND 0.036164f
C595 VPWR.t62 VGND 0.019022f
C596 VPWR.t64 VGND 0.019022f
C597 VPWR.t66 VGND 0.020128f
C598 VPWR.t4 VGND 0.017916f
C599 VPWR.t88 VGND 0.02046f
C600 VPWR.t131 VGND 0.010838f
C601 VPWR.t176 VGND 0.010728f
C602 VPWR.t101 VGND 0.007963f
C603 VPWR.t201 VGND 0.007963f
C604 VPWR.t178 VGND 0.018248f
C605 VPWR.t105 VGND 0.008295f
C606 VPWR.t20 VGND 0.030413f
C607 VPWR.t46 VGND 0.032846f
C608 VPWR.t185 VGND 0.01482f
C609 VPWR.t170 VGND 0.01858f
C610 VPWR.t186 VGND 0.01858f
C611 VPWR.t171 VGND 0.009622f
C612 VPWR.t136 VGND 0.008958f
C613 VPWR.t125 VGND 0.010617f
C614 VPWR.t39 VGND 0.00929f
C615 VPWR.t127 VGND 0.009511f
C616 VPWR.t37 VGND 0.00929f
C617 VPWR.t121 VGND 0.0094f
C618 VPWR.t107 VGND 0.0094f
C619 VPWR.t35 VGND 0.00376f
C620 VPWR.t41 VGND 0.010175f
C621 VPWR.t113 VGND 0.018027f
C622 VPWR.t2 VGND 0.02057f
C623 VPWR.t179 VGND 0.029418f
C624 VPWR.t31 VGND 0.019907f
C625 VPWR.t144 VGND 0.013603f
C626 VPWR.t197 VGND 0.017916f
C627 VPWR.t74 VGND 0.020128f
C628 VPWR.t80 VGND 0.019022f
C629 VPWR.t78 VGND 0.019022f
C630 VPWR.t76 VGND 0.014156f
C631 VPWR.n165 VGND 0.008984f
C632 VPWR.n166 VGND 0.011639f
C633 VPWR.t77 VGND 0.004625f
C634 VPWR.n167 VGND 0.003451f
C635 VPWR.t102 VGND 6.73e-19
C636 VPWR.t132 VGND 0.001016f
C637 VPWR.n168 VGND 0.003036f
C638 VPWR.n169 VGND 0.00455f
C639 VPWR.n170 VGND 0.003133f
C640 VPWR.t67 VGND 0.001485f
C641 VPWR.t5 VGND 0.001094f
C642 VPWR.n171 VGND 0.002785f
C643 VPWR.t208 VGND 0.001485f
C644 VPWR.t150 VGND 0.001094f
C645 VPWR.n172 VGND 0.002785f
C646 VPWR.n173 VGND 0.008976f
C647 VPWR.n174 VGND 0.001201f
C648 VPWR.n175 VGND 0.001157f
C649 VPWR.n176 VGND 0.002063f
C650 VPWR.n178 VGND 0.002063f
C651 VPWR.n179 VGND 0.001728f
C652 VPWR.n180 VGND 9.25e-19
C653 VPWR.n181 VGND 0.001201f
C654 VPWR.n182 VGND 0.001726f
C655 VPWR.t158 VGND 0.002945f
C656 VPWR.t246 VGND 0.006251f
C657 VPWR.n184 VGND 0.016026f
C658 VPWR.t159 VGND 0.002945f
C659 VPWR.n185 VGND 0.008729f
C660 VPWR.t142 VGND 0.002945f
C661 VPWR.t238 VGND 0.006251f
C662 VPWR.n187 VGND 0.016026f
C663 VPWR.t143 VGND 0.002945f
C664 VPWR.n188 VGND 0.008729f
C665 VPWR.n189 VGND 0.007265f
C666 VPWR.t61 VGND 0.004625f
C667 VPWR.n190 VGND 0.003286f
C668 VPWR.n191 VGND 0.004675f
C669 VPWR.t209 VGND 0.004625f
C670 VPWR.n192 VGND 0.009289f
C671 VPWR.n193 VGND 8.04e-19
C672 VPWR.t63 VGND 0.001094f
C673 VPWR.t65 VGND 0.001094f
C674 VPWR.n194 VGND 0.002233f
C675 VPWR.t210 VGND 0.001094f
C676 VPWR.t207 VGND 0.001094f
C677 VPWR.n195 VGND 0.002233f
C678 VPWR.n196 VGND 7.97e-19
C679 VPWR.n197 VGND 0.005139f
C680 VPWR.n198 VGND 0.001201f
C681 VPWR.n199 VGND 9.25e-19
C682 VPWR.n200 VGND 0.001157f
C683 VPWR.n201 VGND 0.001407f
C684 VPWR.n202 VGND 0.001519f
C685 VPWR.n203 VGND 0.001157f
C686 VPWR.n204 VGND 0.00179f
C687 VPWR.n205 VGND 0.002012f
C688 VPWR.n206 VGND 0.105044f
C689 VPWR.n207 VGND 0.002012f
C690 VPWR.n208 VGND 0.00179f
C691 VPWR.n209 VGND 0.001728f
C692 VPWR.n210 VGND 0.002983f
C693 VPWR.n211 VGND 0.002045f
C694 VPWR.n212 VGND 0.001056f
C695 VPWR.n213 VGND 0.001222f
C696 VPWR.t177 VGND 6.73e-19
C697 VPWR.t89 VGND 0.001055f
C698 VPWR.n214 VGND 0.00306f
C699 VPWR.n215 VGND 0.003747f
C700 VPWR.n216 VGND 6.31e-19
C701 VPWR.n217 VGND 0.003451f
C702 VPWR.n218 VGND 0.003451f
C703 VPWR.n219 VGND 8.24e-19
C704 VPWR.n220 VGND 0.001222f
C705 VPWR.n221 VGND 0.00103f
C706 VPWR.n222 VGND 0.002045f
C707 VPWR.n223 VGND 0.001707f
C708 VPWR.n224 VGND 1.53e-19
C709 VPWR.n225 VGND 0.001995f
C710 VPWR.n226 VGND 0.001807f
C711 VPWR.n227 VGND 0.001157f
C712 VPWR.n228 VGND 0.001276f
C713 VPWR.n229 VGND 5.63e-19
C714 VPWR.n230 VGND 0.005361f
C715 VPWR.n231 VGND 0.001434f
C716 VPWR.n232 VGND 0.001201f
C717 VPWR.n233 VGND 0.001276f
C718 VPWR.n234 VGND 0.001157f
C719 VPWR.n235 VGND 9.25e-19
C720 VPWR.n236 VGND 0.002063f
C721 VPWR.n237 VGND 0.001995f
C722 VPWR.n238 VGND 0.001807f
C723 VPWR.n239 VGND 0.001728f
C724 VPWR.n240 VGND 0.001201f
C725 VPWR.n241 VGND 0.002081f
C726 VPWR.n242 VGND 0.003978f
C727 VPWR.n243 VGND 0.004161f
C728 VPWR.n244 VGND 0.00589f
C729 VPWR.n245 VGND 0.0013f
C730 VPWR.n246 VGND 0.003451f
C731 VPWR.n247 VGND 0.002045f
C732 VPWR.n248 VGND 0.003192f
C733 VPWR.n249 VGND 0.004221f
C734 VPWR.n250 VGND 0.003277f
C735 VPWR.t32 VGND 0.002496f
C736 VPWR.t180 VGND 6.07e-19
C737 VPWR.n251 VGND 0.001723f
C738 VPWR.n252 VGND 0.002298f
C739 VPWR.n253 VGND 0.003445f
C740 VPWR.n254 VGND 0.003627f
C741 VPWR.n255 VGND 0.003451f
C742 VPWR.n256 VGND 0.003451f
C743 VPWR.n257 VGND 0.003433f
C744 VPWR.n258 VGND 0.004216f
C745 VPWR.n259 VGND 0.002222f
C746 VPWR.n260 VGND 0.004464f
C747 VPWR.t42 VGND 0.004625f
C748 VPWR.n261 VGND 0.0055f
C749 VPWR.n262 VGND 0.001407f
C750 VPWR.n263 VGND 0.001157f
C751 VPWR.n264 VGND 0.002063f
C752 VPWR.n265 VGND 9.25e-19
C753 VPWR.t108 VGND 0.001055f
C754 VPWR.t122 VGND 0.001055f
C755 VPWR.n266 VGND 0.002317f
C756 VPWR.n267 VGND 0.003114f
C757 VPWR.t36 VGND 0.001094f
C758 VPWR.t38 VGND 0.001094f
C759 VPWR.n268 VGND 0.00223f
C760 VPWR.t128 VGND 0.001055f
C761 VPWR.t126 VGND 0.001055f
C762 VPWR.n269 VGND 0.00227f
C763 VPWR.n270 VGND 0.003538f
C764 VPWR.n271 VGND 0.002045f
C765 VPWR.t40 VGND 0.001485f
C766 VPWR.t137 VGND 0.001094f
C767 VPWR.n272 VGND 0.002741f
C768 VPWR.n273 VGND 0.003861f
C769 VPWR.t47 VGND 0.002921f
C770 VPWR.n274 VGND 0.005145f
C771 VPWR.n275 VGND 0.001728f
C772 VPWR.t239 VGND 0.017175f
C773 VPWR.n276 VGND 0.00906f
C774 VPWR.n277 VGND 0.001201f
C775 VPWR.n278 VGND 0.001807f
C776 VPWR.n279 VGND 0.001157f
C777 VPWR.n280 VGND 0.002063f
C778 VPWR.n282 VGND 0.002012f
C779 VPWR.n283 VGND 0.002063f
C780 VPWR.n284 VGND 0.001157f
C781 VPWR.n285 VGND 0.001201f
C782 VPWR.t152 VGND -1.44e-20
C783 VPWR.t100 VGND 9e-19
C784 VPWR.n286 VGND 0.003971f
C785 VPWR.t154 VGND 0.004284f
C786 VPWR.n287 VGND 0.006081f
C787 VPWR.n288 VGND 0.001726f
C788 VPWR.n289 VGND 0.001501f
C789 VPWR.n290 VGND 0.003451f
C790 VPWR.n291 VGND 0.00435f
C791 VPWR.n292 VGND 0.003451f
C792 VPWR.n293 VGND 0.003192f
C793 VPWR.n294 VGND 0.001332f
C794 VPWR.n295 VGND 0.001157f
C795 VPWR.n296 VGND 0.002063f
C796 VPWR.n297 VGND 0.002063f
C797 VPWR.n298 VGND 0.001728f
C798 VPWR.n299 VGND 9.25e-19
C799 VPWR.n300 VGND 0.001201f
C800 VPWR.n301 VGND 9.25e-19
C801 VPWR.n302 VGND 0.001157f
C802 VPWR.n303 VGND 0.001726f
C803 VPWR.n304 VGND 0.003395f
C804 VPWR.t243 VGND 0.012191f
C805 VPWR.n305 VGND 9.52e-19
C806 VPWR.n306 VGND 0.001728f
C807 VPWR.t163 VGND 0.004284f
C808 VPWR.t212 VGND 9e-19
C809 VPWR.t161 VGND -1.44e-20
C810 VPWR.n307 VGND 0.003971f
C811 VPWR.n308 VGND 0.005383f
C812 VPWR.n309 VGND 0.001201f
C813 VPWR.n310 VGND 9.25e-19
C814 VPWR.n311 VGND 9.25e-19
C815 VPWR.n312 VGND 4.53e-19
C816 VPWR.n313 VGND 0.001157f
C817 VPWR.n314 VGND 0.001407f
C818 VPWR.n315 VGND 0.001669f
C819 VPWR.t71 VGND 0.022015f
C820 VPWR.t26 VGND 0.024148f
C821 VPWR.t133 VGND 0.013987f
C822 VPWR.t111 VGND 0.010663f
C823 VPWR.t135 VGND 0.016559f
C824 VPWR.t166 VGND 0.016057f
C825 VPWR.t138 VGND 0.017311f
C826 VPWR.t99 VGND 0.010035f
C827 VPWR.t151 VGND 0.011227f
C828 VPWR.t153 VGND 0.013046f
C829 VPWR.t155 VGND 0.069244f
C830 VPWR.t94 VGND 0.023207f
C831 VPWR.t162 VGND 0.015053f
C832 VPWR.t160 VGND 0.011227f
C833 VPWR.t211 VGND 0.007903f
C834 VPWR.n316 VGND 0.013384f
C835 VPWR.n317 VGND 0.001036f
C836 VPWR.n318 VGND 0.003451f
C837 VPWR.t167 VGND 0.001803f
C838 VPWR.n319 VGND 0.001016f
C839 VPWR.n320 VGND 0.001728f
C840 VPWR.t112 VGND 6.73e-19
C841 VPWR.t134 VGND 0.001055f
C842 VPWR.n321 VGND 0.003104f
C843 VPWR.t228 VGND 0.006139f
C844 VPWR.n322 VGND 0.009289f
C845 VPWR.n323 VGND 0.007632f
C846 VPWR.t28 VGND 0.002945f
C847 VPWR.n324 VGND 0.005121f
C848 VPWR.n325 VGND 0.003462f
C849 VPWR.n326 VGND 9.25e-19
C850 VPWR.n327 VGND 0.001519f
C851 VPWR.n328 VGND 5.25e-19
C852 VPWR.n329 VGND 0.001407f
C853 VPWR.n330 VGND 0.001157f
C854 VPWR.n331 VGND 0.002063f
C855 VPWR.n332 VGND 9.25e-19
C856 VPWR.n333 VGND 0.001807f
C857 VPWR.n334 VGND 0.001157f
C858 VPWR.n335 VGND 0.001407f
C859 VPWR.n336 VGND 0.001201f
C860 VPWR.n337 VGND 9.72e-19
C861 VPWR.n338 VGND 0.004899f
C862 VPWR.n339 VGND 0.002983f
C863 VPWR.n340 VGND 0.003451f
C864 VPWR.n341 VGND 0.003451f
C865 VPWR.n342 VGND 0.001222f
C866 VPWR.n343 VGND 0.00107f
C867 VPWR.n344 VGND 0.006009f
C868 VPWR.n345 VGND 0.002026f
C869 VPWR.n346 VGND 0.003151f
C870 VPWR.n347 VGND 0.002195f
C871 VPWR.n348 VGND 0.00103f
C872 VPWR.n349 VGND 0.007308f
C873 VPWR.n350 VGND 8.57e-19
C874 VPWR.n351 VGND 4.31e-19
C875 VPWR.n352 VGND 0.001276f
C876 VPWR.n353 VGND 0.001157f
C877 VPWR.n354 VGND 0.001807f
C878 VPWR.n355 VGND 0.001995f
C879 VPWR.n356 VGND 0.002063f
C880 VPWR.n357 VGND 0.002063f
C881 VPWR.n358 VGND 0.001995f
C882 VPWR.n359 VGND 0.001807f
C883 VPWR.n360 VGND 0.001157f
C884 VPWR.n361 VGND 0.001726f
C885 VPWR.n362 VGND 0.001201f
C886 VPWR.n363 VGND 7.97e-19
C887 VPWR.n364 VGND 0.0061f
C888 VPWR.n365 VGND 0.003414f
C889 VPWR.n366 VGND 0.002176f
C890 VPWR.n367 VGND 0.003001f
C891 VPWR.n368 VGND 0.003462f
C892 VPWR.t95 VGND 0.002921f
C893 VPWR.n369 VGND 0.00288f
C894 VPWR.n370 VGND 0.011027f
C895 VPWR.n371 VGND 0.006795f
C896 VPWR.t96 VGND 0.002921f
C897 VPWR.n372 VGND 0.005145f
C898 VPWR.n373 VGND 0.008765f
C899 VPWR.n374 VGND 0.003451f
C900 VPWR.n375 VGND 0.002045f
C901 VPWR.n376 VGND 0.003114f
C902 VPWR.n377 VGND 0.001687f
C903 VPWR.t156 VGND 0.003214f
C904 VPWR.n378 VGND 0.002497f
C905 VPWR.n379 VGND 0.004208f
C906 VPWR.t245 VGND 0.04257f
C907 VPWR.n380 VGND 0.019884f
C908 VPWR.n381 VGND 0.001201f
C909 VPWR.n382 VGND 0.003333f
C910 VPWR.n383 VGND 0.00435f
C911 VPWR.n384 VGND 0.001201f
C912 VPWR.n385 VGND 0.001726f
C913 VPWR.n386 VGND 0.001157f
C914 VPWR.n387 VGND 0.001807f
C915 VPWR.n388 VGND 0.001995f
C916 VPWR.n389 VGND 0.074031f
C917 VPWR.n390 VGND 0.001995f
C918 VPWR.n391 VGND 0.001807f
C919 VPWR.n392 VGND 0.001597f
C920 VPWR.n393 VGND 0.00212f
C921 VPWR.n394 VGND 0.003451f
C922 VPWR.n395 VGND 0.00435f
C923 VPWR.n396 VGND 0.00435f
C924 VPWR.n397 VGND 0.00435f
C925 VPWR.n398 VGND 0.003451f
C926 VPWR.n399 VGND 0.003451f
C927 VPWR.n400 VGND 0.003451f
C928 VPWR.n401 VGND 0.00435f
C929 VPWR.n402 VGND 0.004208f
C930 VPWR.t157 VGND 0.003214f
C931 VPWR.n403 VGND 0.002497f
C932 VPWR.n404 VGND 0.001572f
C933 VPWR.n405 VGND 0.002045f
C934 VPWR.n406 VGND 0.001201f
C935 VPWR.n407 VGND 0.001409f
C936 VPWR.n408 VGND 0.00179f
C937 VPWR.n409 VGND 0.001157f
C938 VPWR.n410 VGND 0.002063f
C939 VPWR.n411 VGND 9.25e-19
C940 VPWR.n412 VGND 9.25e-19
C941 VPWR.n413 VGND 0.001157f
C942 VPWR.n414 VGND 0.001426f
C943 VPWR.n415 VGND 0.001201f
C944 VPWR.n416 VGND 7.97e-19
C945 VPWR.n417 VGND 0.005383f
C946 VPWR.t139 VGND 0.002945f
C947 VPWR.n418 VGND 0.001723f
C948 VPWR.n419 VGND 0.002137f
C949 VPWR.t234 VGND 0.006139f
C950 VPWR.n420 VGND 0.009289f
C951 VPWR.t140 VGND 0.002945f
C952 VPWR.n421 VGND 0.007954f
C953 VPWR.n422 VGND 0.007632f
C954 VPWR.n423 VGND 0.003451f
C955 VPWR.n424 VGND 0.003133f
C956 VPWR.n425 VGND 0.003462f
C957 VPWR.n426 VGND 9.65e-19
C958 VPWR.n427 VGND 0.001144f
C959 VPWR.n428 VGND 0.001728f
C960 VPWR.n429 VGND 0.00179f
C961 VPWR.n430 VGND 0.002012f
C962 VPWR.n431 VGND 0.074031f
C963 VPWR.n432 VGND 0.001995f
C964 VPWR.n433 VGND 0.002063f
C965 VPWR.n434 VGND 0.001728f
C966 VPWR.n435 VGND 9.25e-19
C967 VPWR.n436 VGND 0.001201f
C968 VPWR.n437 VGND 0.001426f
C969 VPWR.n438 VGND 0.007478f
C970 VPWR.n439 VGND 0.003451f
C971 VPWR.t241 VGND 0.04257f
C972 VPWR.t224 VGND 0.04257f
C973 VPWR.n440 VGND 0.007478f
C974 VPWR.n441 VGND 0.00212f
C975 VPWR.t214 VGND 0.003214f
C976 VPWR.t70 VGND 0.003214f
C977 VPWR.n442 VGND 0.004383f
C978 VPWR.n443 VGND 0.001726f
C979 VPWR.n444 VGND 9.25e-19
C980 VPWR.n445 VGND 0.001409f
C981 VPWR.n446 VGND 0.002012f
C982 VPWR.n447 VGND 0.00179f
C983 VPWR.n448 VGND 0.001201f
C984 VPWR.n449 VGND 0.007478f
C985 VPWR.n450 VGND 0.003451f
C986 VPWR.t236 VGND 0.04257f
C987 VPWR.t222 VGND 0.04257f
C988 VPWR.n451 VGND 0.039157f
C989 VPWR.n452 VGND 0.003414f
C990 VPWR.n453 VGND 0.007234f
C991 VPWR.n454 VGND 0.007478f
C992 VPWR.n455 VGND 0.005731f
C993 VPWR.n456 VGND 0.003451f
C994 VPWR.n457 VGND 0.003451f
C995 VPWR.n458 VGND 0.005487f
C996 VPWR.n459 VGND 0.007478f
C997 VPWR.n460 VGND 0.007478f
C998 VPWR.n461 VGND 0.003451f
C999 VPWR.n462 VGND 0.003451f
C1000 VPWR.n463 VGND 0.001728f
C1001 VPWR.n464 VGND 0.003433f
C1002 VPWR.n465 VGND 0.007478f
C1003 VPWR.n466 VGND 0.007478f
C1004 VPWR.n467 VGND 0.007234f
C1005 VPWR.n468 VGND 0.001201f
C1006 VPWR.n469 VGND 0.001726f
C1007 VPWR.n470 VGND 0.001157f
C1008 VPWR.n471 VGND 0.001157f
C1009 VPWR.n472 VGND 9.25e-19
C1010 VPWR.n473 VGND 0.002063f
C1011 VPWR.n475 VGND 0.002063f
C1012 VPWR.n476 VGND 0.002012f
C1013 VPWR.n477 VGND 0.00179f
C1014 VPWR.n478 VGND 0.001157f
C1015 VPWR.n479 VGND 3.19e-19
C1016 VPWR.n480 VGND 0.001201f
C1017 VPWR.n481 VGND 0.002824f
C1018 VPWR.n482 VGND 0.002762f
C1019 VPWR.t92 VGND 0.003214f
C1020 VPWR.t86 VGND 0.003214f
C1021 VPWR.n483 VGND 0.004383f
C1022 VPWR.n484 VGND 0.007234f
C1023 VPWR.n485 VGND 0.003451f
C1024 VPWR.n486 VGND 0.003451f
C1025 VPWR.n487 VGND 0.003451f
C1026 VPWR.n488 VGND 0.005731f
C1027 VPWR.n489 VGND 0.039157f
C1028 VPWR.n490 VGND 0.005487f
C1029 VPWR.n491 VGND 0.007478f
C1030 VPWR.n492 VGND 0.003451f
C1031 VPWR.n493 VGND 0.003451f
C1032 VPWR.n494 VGND 0.003001f
C1033 VPWR.n495 VGND 0.007478f
C1034 VPWR.n496 VGND 0.007478f
C1035 VPWR.t93 VGND 0.003214f
C1036 VPWR.t87 VGND 0.003214f
C1037 VPWR.n497 VGND 0.004383f
C1038 VPWR.n498 VGND 0.001501f
C1039 VPWR.t44 VGND 0.002945f
C1040 VPWR.t244 VGND 0.006251f
C1041 VPWR.n500 VGND 0.016026f
C1042 VPWR.t45 VGND 0.002945f
C1043 VPWR.n501 VGND 0.008729f
C1044 VPWR.t52 VGND 0.002945f
C1045 VPWR.t227 VGND 0.006251f
C1046 VPWR.n503 VGND 0.016026f
C1047 VPWR.t53 VGND 0.002945f
C1048 VPWR.n504 VGND 0.008729f
C1049 VPWR.n505 VGND 0.00358f
C1050 VPWR.n506 VGND 0.007359f
C1051 VPWR.n507 VGND 0.002655f
C1052 VPWR.n508 VGND 0.001144f
C1053 VPWR.n509 VGND 0.001157f
C1054 VPWR.n510 VGND 0.002063f
C1055 VPWR.n511 VGND 9.25e-19
C1056 VPWR.n512 VGND 0.001157f
C1057 VPWR.n513 VGND 0.001807f
C1058 VPWR.n514 VGND 0.001728f
C1059 VPWR.n515 VGND 0.001201f
C1060 VPWR.n516 VGND 0.007234f
C1061 VPWR.n517 VGND 0.007478f
C1062 VPWR.n518 VGND 0.001201f
C1063 VPWR.n519 VGND 0.001726f
C1064 VPWR.n520 VGND 0.001157f
C1065 VPWR.n521 VGND 0.001807f
C1066 VPWR.n522 VGND 0.001995f
C1067 VPWR.n523 VGND 0.136057f
C1068 VPWR.n524 VGND 0.001995f
C1069 VPWR.n525 VGND 0.002063f
C1070 VPWR.n526 VGND 0.001728f
C1071 VPWR.n527 VGND 9.25e-19
C1072 VPWR.n528 VGND 0.001201f
C1073 VPWR.n529 VGND 0.001426f
C1074 VPWR.n530 VGND 0.003277f
C1075 VPWR.n531 VGND 0.003133f
C1076 VPWR.t149 VGND 0.003214f
C1077 VPWR.n532 VGND 0.002069f
C1078 VPWR.n533 VGND 0.003451f
C1079 VPWR.t50 VGND 0.003214f
C1080 VPWR.n534 VGND 0.004061f
C1081 VPWR.n535 VGND 0.001409f
C1082 VPWR.t217 VGND 0.003214f
C1083 VPWR.n536 VGND 0.004061f
C1084 VPWR.n537 VGND 0.001726f
C1085 VPWR.n538 VGND 0.005487f
C1086 VPWR.n539 VGND 0.007234f
C1087 VPWR.n540 VGND 0.001201f
C1088 VPWR.n541 VGND 0.001726f
C1089 VPWR.n542 VGND 9.25e-19
C1090 VPWR.n543 VGND 0.001157f
C1091 VPWR.n544 VGND 0.002063f
C1092 VPWR.n545 VGND 9.25e-19
C1093 VPWR.n546 VGND 0.001807f
C1094 VPWR.n547 VGND 0.001157f
C1095 VPWR.n548 VGND 3.19e-19
C1096 VPWR.n549 VGND 0.001201f
C1097 VPWR.n550 VGND 0.003402f
C1098 VPWR.n551 VGND 0.003374f
C1099 VPWR.n552 VGND 0.00212f
C1100 VPWR.n553 VGND 0.003451f
C1101 VPWR.n554 VGND 0.007234f
C1102 VPWR.n555 VGND 0.007478f
C1103 VPWR.t231 VGND 0.04257f
C1104 VPWR.n556 VGND 0.021204f
C1105 VPWR.n557 VGND 0.005731f
C1106 VPWR.n558 VGND 0.003451f
C1107 VPWR.n559 VGND 0.002045f
C1108 VPWR.n560 VGND 0.003527f
C1109 VPWR.n561 VGND 0.004099f
C1110 VPWR.t200 VGND 0.002496f
C1111 VPWR.t116 VGND 6.07e-19
C1112 VPWR.n562 VGND 0.001723f
C1113 VPWR.n563 VGND 0.002298f
C1114 VPWR.n564 VGND 0.003445f
C1115 VPWR.n565 VGND 0.003627f
C1116 VPWR.n566 VGND 0.003451f
C1117 VPWR.n567 VGND 0.003001f
C1118 VPWR.n568 VGND 0.003647f
C1119 VPWR.n569 VGND 0.004216f
C1120 VPWR.t1 VGND 6.73e-19
C1121 VPWR.t169 VGND 4.43e-19
C1122 VPWR.n570 VGND 0.001149f
C1123 VPWR.t51 VGND 0.003214f
C1124 VPWR.n571 VGND 0.002497f
C1125 VPWR.n572 VGND 0.001501f
C1126 VPWR.t29 VGND 0.002945f
C1127 VPWR.t233 VGND 0.006251f
C1128 VPWR.n574 VGND 0.016026f
C1129 VPWR.t30 VGND 0.002945f
C1130 VPWR.n575 VGND 0.008729f
C1131 VPWR.t7 VGND 0.002945f
C1132 VPWR.t220 VGND 0.006251f
C1133 VPWR.n577 VGND 0.016026f
C1134 VPWR.t8 VGND 0.002945f
C1135 VPWR.n578 VGND 0.008729f
C1136 VPWR.n579 VGND 0.003421f
C1137 VPWR.n580 VGND 0.007364f
C1138 VPWR.n581 VGND 0.001562f
C1139 VPWR.n582 VGND 0.001144f
C1140 VPWR.n583 VGND 0.001157f
C1141 VPWR.n584 VGND 0.002063f
C1142 VPWR.n585 VGND 9.25e-19
C1143 VPWR.n586 VGND 0.001157f
C1144 VPWR.n587 VGND 0.001807f
C1145 VPWR.n588 VGND 0.001409f
C1146 VPWR.n589 VGND 6.19e-19
C1147 VPWR.n590 VGND 0.004161f
C1148 VPWR.n591 VGND 0.004464f
C1149 VPWR.n592 VGND 0.002222f
C1150 VPWR.n593 VGND 0.001201f
C1151 VPWR.n594 VGND 0.001726f
C1152 VPWR.n595 VGND 0.001157f
C1153 VPWR.n596 VGND 0.001807f
C1154 VPWR.n597 VGND 0.001995f
C1155 VPWR.n598 VGND 0.136057f
C1156 VPWR.n599 VGND 9.25e-19
C1157 VPWR.n600 VGND 0.001157f
C1158 VPWR.n601 VGND 0.001426f
C1159 VPWR.n602 VGND 0.001501f
C1160 VPWR.n603 VGND 0.001201f
C1161 VPWR.n604 VGND 0.008765f
C1162 VPWR.t48 VGND 0.002921f
C1163 VPWR.n605 VGND 0.005145f
C1164 VPWR.t202 VGND 0.002945f
C1165 VPWR.t219 VGND 0.006251f
C1166 VPWR.n607 VGND 0.016026f
C1167 VPWR.t203 VGND 0.002945f
C1168 VPWR.n608 VGND 0.008729f
C1169 VPWR.t21 VGND 0.002945f
C1170 VPWR.t242 VGND 0.006251f
C1171 VPWR.n610 VGND 0.016026f
C1172 VPWR.t22 VGND 0.002945f
C1173 VPWR.n611 VGND 0.008729f
C1174 VPWR.n612 VGND 0.003398f
C1175 VPWR.n613 VGND 0.007358f
C1176 VPWR.n614 VGND 0.003207f
C1177 VPWR.n615 VGND 0.001144f
C1178 VPWR.n616 VGND 0.001728f
C1179 VPWR.n617 VGND 0.001807f
C1180 VPWR.n618 VGND 0.001995f
C1181 VPWR.n619 VGND 0.105044f
C1182 VPWR.n620 VGND 0.001995f
C1183 VPWR.n621 VGND 0.002063f
C1184 VPWR.n622 VGND 9.25e-19
C1185 VPWR.n623 VGND 0.001157f
C1186 VPWR.n624 VGND 0.001726f
C1187 VPWR.n625 VGND 0.001201f
C1188 VPWR.n626 VGND 0.00906f
C1189 VPWR.n627 VGND 0.023314f
C1190 VPWR.n628 VGND 0.003001f
C1191 VPWR.n629 VGND 0.003133f
C1192 VPWR.n630 VGND 0.003462f
C1193 VPWR.n631 VGND 0.001138f
C1194 VPWR.n632 VGND 6.51e-19
C1195 VPWR.n633 VGND 0.003451f
C1196 VPWR.n634 VGND 0.003451f
C1197 VPWR.n635 VGND 8.44e-19
C1198 VPWR.n636 VGND 0.007373f
C1199 VPWR.n637 VGND 7.57e-19
C1200 VPWR.n638 VGND 0.001594f
C1201 VPWR.n639 VGND 8.63e-19
C1202 VPWR.n640 VGND 0.001409f
C1203 VPWR.n641 VGND 0.001807f
C1204 VPWR.n642 VGND 0.001157f
C1205 VPWR.n643 VGND 3.19e-19
C1206 VPWR.n644 VGND 0.001201f
C1207 VPWR.n645 VGND 0.001661f
C1208 VPWR.t146 VGND 0.003214f
C1209 VPWR.n646 VGND 0.002497f
C1210 VPWR.n647 VGND 0.004161f
C1211 VPWR.n648 VGND 8.63e-19
C1212 VPWR.n649 VGND 0.001726f
C1213 VPWR.n650 VGND 0.001157f
C1214 VPWR.n651 VGND 0.001807f
C1215 VPWR.n652 VGND 0.001995f
C1216 VPWR.n653 VGND 0.105044f
C1217 VPWR.n654 VGND 0.136057f
C1218 VPWR.n655 VGND 0.001995f
C1219 VPWR.n656 VGND 0.001807f
C1220 VPWR.n657 VGND 0.001728f
C1221 VPWR.n658 VGND 0.003433f
C1222 VPWR.n659 VGND 0.005731f
C1223 VPWR.n660 VGND 0.007478f
C1224 VPWR.n661 VGND 0.007234f
C1225 VPWR.n662 VGND 0.003451f
C1226 VPWR.n663 VGND 0.003133f
C1227 VPWR.n664 VGND 0.002045f
C1228 VPWR.n665 VGND 0.005124f
C1229 VPWR.t59 VGND 0.002921f
C1230 VPWR.n666 VGND 0.003463f
C1231 VPWR.n667 VGND 0.023405f
C1232 VPWR.n668 VGND 0.009339f
C1233 VPWR.n669 VGND 0.012188f
C1234 VPWR.n670 VGND 0.003414f
C1235 VPWR.n671 VGND 0.001728f
C1236 VPWR.n672 VGND 0.00179f
C1237 VPWR.n673 VGND 0.002012f
C1238 VPWR.n674 VGND 0.136057f
C1239 VPWR.n675 VGND 0.002063f
C1240 VPWR.n676 VGND 0.001157f
C1241 VPWR.n677 VGND 9.25e-19
C1242 VPWR.n678 VGND 0.001276f
C1243 VPWR.n679 VGND 0.001157f
C1244 VPWR.n680 VGND 0.001807f
C1245 VPWR.n681 VGND 0.001995f
C1246 VPWR.n682 VGND 0.136057f
C1247 VPWR.n683 VGND 0.001995f
C1248 VPWR.n684 VGND 0.001807f
C1249 VPWR.n685 VGND 0.001157f
C1250 VPWR.n686 VGND 0.001726f
C1251 VPWR.n687 VGND 0.001201f
C1252 VPWR.n688 VGND 0.002594f
C1253 VPWR.n689 VGND 0.01089f
C1254 VPWR.n690 VGND 0.00182f
C1255 VPWR.n691 VGND 0.002513f
C1256 VPWR.n692 VGND 0.005097f
C1257 VPWR.t206 VGND 0.002965f
C1258 VPWR.n693 VGND 0.002875f
C1259 VPWR.n694 VGND 0.012269f
C1260 VPWR.t221 VGND 0.012354f
C1261 VPWR.n695 VGND 0.013501f
C1262 VPWR.t205 VGND 0.002921f
C1263 VPWR.n696 VGND 0.004241f
C1264 VPWR.n697 VGND 0.008762f
C1265 VPWR.n698 VGND 0.002311f
C1266 VPWR.n699 VGND 0.001857f
C1267 VPWR.n700 VGND 6.78e-19
C1268 VPWR.n701 VGND 0.00105f
C1269 VPWR.n702 VGND 0.002045f
C1270 VPWR.n703 VGND 0.002983f
C1271 VPWR.n704 VGND 2.13e-19
C1272 VPWR.n705 VGND 0.004326f
C1273 VPWR.n706 VGND 9.04e-19
C1274 VPWR.n707 VGND 0.001201f
C1275 VPWR.n708 VGND 0.001726f
C1276 VPWR.n709 VGND 0.001157f
C1277 VPWR.n710 VGND 0.002063f
C1278 VPWR.n711 VGND 9.25e-19
C1279 VPWR.n712 VGND 0.001157f
C1280 VPWR.n713 VGND 0.001407f
C1281 VPWR.n714 VGND 0.001519f
C1282 VPWR.n715 VGND 0.001157f
C1283 VPWR.n716 VGND 0.001807f
C1284 VPWR.n717 VGND 0.001995f
C1285 VPWR.n718 VGND 0.136057f
C1286 VPWR.n719 VGND 0.074031f
C1287 VPWR.n720 VGND 0.001995f
C1288 VPWR.n721 VGND 0.001807f
C1289 VPWR.n722 VGND 0.001728f
C1290 VPWR.n723 VGND 0.00257f
C1291 VPWR.n724 VGND 0.003377f
C1292 VPWR.n725 VGND 0.003377f
C1293 VPWR.t73 VGND 0.002945f
C1294 VPWR.n726 VGND 0.001723f
C1295 VPWR.n727 VGND 0.009289f
C1296 VPWR.n728 VGND 0.007632f
C1297 VPWR.n729 VGND 0.003133f
.ends

